library verilog;
use verilog.vl_types.all;
entity t_alu is
end t_alu;
