library verilog;
use verilog.vl_types.all;
entity t_Add_4bitRCA is
end t_Add_4bitRCA;
