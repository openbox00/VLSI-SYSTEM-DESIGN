library verilog;
use verilog.vl_types.all;
entity INST_MEM is
    generic(
        IM_SIZE         : integer := 104857600
    );
    port(
        clk             : in     vl_logic;
        pc              : in     vl_logic_vector(31 downto 0);
        inst_out        : out    vl_logic_vector(31 downto 0)
    );
end INST_MEM;
