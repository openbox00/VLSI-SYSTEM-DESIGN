`timescale 1ns/10ps
module ALU_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [1:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] , n1,
         n2, n3, n4;

  MX2X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S0(n2), .Y(\ML_int[1][22] ) );
  MX2X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S0(n2), .Y(\ML_int[1][24] ) );
  MX2X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S0(n2), .Y(\ML_int[1][25] ) );
  MX2X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S0(n2), .Y(\ML_int[1][26] ) );
  MX2X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S0(n2), .Y(\ML_int[1][23] ) );
  MX2X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S0(n2), .Y(\ML_int[1][27] ) );
  MX2X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S0(n2), .Y(\ML_int[1][28] ) );
  MX2X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S0(n2), .Y(\ML_int[1][29] ) );
  MX2X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S0(n2), .Y(\ML_int[1][31] ) );
  MX2X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S0(SH[1]), .Y(
        B[31]) );
  MX2X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S0(n2), .Y(\ML_int[1][15] ) );
  MX2X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S0(n2), .Y(\ML_int[1][16] ) );
  MX2X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S0(n2), .Y(\ML_int[1][12] ) );
  MX2X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S0(n2), .Y(\ML_int[1][18] ) );
  MX2X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S0(n2), .Y(\ML_int[1][14] ) );
  MX2X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S0(n2), .Y(\ML_int[1][21] ) );
  MX2X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S0(n2), .Y(\ML_int[1][20] ) );
  MX2X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S0(n2), .Y(\ML_int[1][13] ) );
  MX2X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S0(n2), .Y(\ML_int[1][17] ) );
  MX2X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S0(n2), .Y(\ML_int[1][19] ) );
  MX2X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S0(n1), .Y(\ML_int[1][1] ) );
  MX2X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S0(n2), .Y(\ML_int[1][30] ) );
  MX2X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S0(SH[1]), .Y(
        B[30]) );
  MX2X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S0(SH[1]), .Y(
        B[29]) );
  MX2X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S0(SH[1]), .Y(
        B[28]) );
  MX2X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S0(SH[1]), .Y(
        B[27]) );
  MX2X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S0(SH[1]), .Y(
        B[26]) );
  MX2X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S0(SH[1]), .Y(
        B[25]) );
  MX2X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S0(SH[1]), .Y(
        B[24]) );
  MX2X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S0(SH[1]), .Y(
        B[23]) );
  MX2X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S0(SH[1]), .Y(
        B[22]) );
  MX2X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S0(SH[1]), .Y(
        B[21]) );
  MX2X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S0(SH[1]), .Y(
        B[20]) );
  MX2X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S0(SH[1]), .Y(
        B[19]) );
  MX2X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S0(SH[1]), .Y(
        B[18]) );
  MX2X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S0(SH[1]), .Y(
        B[17]) );
  MX2X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S0(SH[1]), .Y(
        B[16]) );
  MX2X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S0(SH[1]), .Y(
        B[15]) );
  MX2X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S0(SH[1]), .Y(
        B[14]) );
  MX2X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S0(SH[1]), .Y(
        B[13]) );
  MX2X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S0(SH[1]), .Y(
        B[12]) );
  MX2X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S0(SH[1]), .Y(
        B[11]) );
  MX2X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S0(SH[1]), .Y(
        B[10]) );
  MX2X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S0(SH[1]), .Y(B[9])
         );
  MX2X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S0(SH[1]), .Y(B[8])
         );
  MX2X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S0(SH[1]), .Y(B[7])
         );
  MX2X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S0(SH[1]), .Y(B[6])
         );
  MX2X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S0(SH[1]), .Y(B[5])
         );
  MX2X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S0(SH[1]), .Y(B[4])
         );
  MX2X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S0(SH[1]), .Y(B[3])
         );
  MX2X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S0(SH[1]), .Y(B[2])
         );
  MX2X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S0(n1), .Y(\ML_int[1][2] ) );
  MX2X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S0(n2), .Y(\ML_int[1][4] ) );
  MX2X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S0(n1), .Y(\ML_int[1][3] ) );
  MX2X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S0(n2), .Y(\ML_int[1][5] ) );
  MX2X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S0(n2), .Y(\ML_int[1][6] ) );
  MX2X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S0(n2), .Y(\ML_int[1][11] ) );
  MX2X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S0(SH[0]), .Y(\ML_int[1][7] ) );
  MX2X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S0(SH[0]), .Y(\ML_int[1][8] ) );
  MX2X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S0(SH[0]), .Y(\ML_int[1][9] ) );
  MX2X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S0(n2), .Y(\ML_int[1][10] ) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n2) );
  INVX1 U5 ( .A(SH[0]), .Y(n3) );
  NOR2BX1 U6 ( .AN(\ML_int[1][1] ), .B(SH[1]), .Y(B[1]) );
  NOR2X1 U7 ( .A(SH[1]), .B(n4), .Y(B[0]) );
  INVX1 U8 ( .A(n4), .Y(\ML_int[1][0] ) );
  NAND2X1 U9 ( .A(A[0]), .B(n3), .Y(n4) );
endmodule


module ALU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] ;

  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        SUM[5]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        SUM[6]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        SUM[7]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        SUM[8]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(\carry[31] ), .Y(SUM[31]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(\carry[1] ) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module ALU_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] , \B_not[31] , \B_not[30] , \B_not[29] , \B_not[28] ,
         \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] , \B_not[23] ,
         \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] , \B_not[18] ,
         \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] , \B_not[13] ,
         \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] , \B_not[8] ,
         \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] , \B_not[3] ,
         \B_not[2] , \B_not[1] , \B_not[0] ;

  ADDFX2 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), 
        .S(DIFF[5]) );
  ADDFX2 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), 
        .S(DIFF[3]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), 
        .S(DIFF[1]) );
  ADDFX2 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), 
        .S(DIFF[2]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(\B_not[4] ), .CI(\carry[4] ), .CO(\carry[5] ), 
        .S(DIFF[4]) );
  ADDFX2 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), .S(DIFF[14]) );
  ADDFX2 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), .S(DIFF[15]) );
  ADDFX2 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), .S(DIFF[17]) );
  ADDFX2 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), .S(DIFF[11]) );
  ADDFX2 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), .S(DIFF[20]) );
  ADDFX2 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), .S(DIFF[19]) );
  ADDFX2 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), .S(DIFF[13]) );
  ADDFX2 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), .S(DIFF[21]) );
  ADDFX2 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), .S(DIFF[12]) );
  ADDFX2 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), .S(DIFF[18]) );
  ADDFX2 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), .S(DIFF[16]) );
  ADDFX2 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), .S(DIFF[10]) );
  ADDFX2 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), .S(DIFF[23]) );
  ADDFX2 U2_30 ( .A(A[30]), .B(\B_not[30] ), .CI(\carry[30] ), .CO(\carry[31] ), .S(DIFF[30]) );
  ADDFX2 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), .S(DIFF[24]) );
  ADDFX2 U2_29 ( .A(A[29]), .B(\B_not[29] ), .CI(\carry[29] ), .CO(\carry[30] ), .S(DIFF[29]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), 
        .S(DIFF[6]) );
  ADDFX2 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), .S(DIFF[25]) );
  ADDFX2 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), .S(DIFF[22]) );
  ADDFX2 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), .S(DIFF[27]) );
  ADDFX2 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), .S(DIFF[26]) );
  ADDFX2 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), .S(DIFF[28]) );
  ADDFX2 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), 
        .S(DIFF[7]) );
  ADDFX2 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), 
        .S(DIFF[8]) );
  ADDFX2 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  XOR3X2 U2_31 ( .A(A[31]), .B(\B_not[31] ), .C(\carry[31] ), .Y(DIFF[31]) );
  OR2X1 U1 ( .A(\B_not[0] ), .B(A[0]), .Y(\carry[1] ) );
  XNOR2X1 U2 ( .A(A[0]), .B(\B_not[0] ), .Y(DIFF[0]) );
  INVX1 U3 ( .A(B[9]), .Y(\B_not[9] ) );
  INVX1 U4 ( .A(B[8]), .Y(\B_not[8] ) );
  INVX1 U5 ( .A(B[7]), .Y(\B_not[7] ) );
  INVX1 U6 ( .A(B[6]), .Y(\B_not[6] ) );
  INVX1 U7 ( .A(B[5]), .Y(\B_not[5] ) );
  INVX1 U8 ( .A(B[4]), .Y(\B_not[4] ) );
  INVX1 U9 ( .A(B[3]), .Y(\B_not[3] ) );
  INVX1 U10 ( .A(B[31]), .Y(\B_not[31] ) );
  INVX1 U11 ( .A(B[30]), .Y(\B_not[30] ) );
  INVX1 U12 ( .A(B[2]), .Y(\B_not[2] ) );
  INVX1 U13 ( .A(B[29]), .Y(\B_not[29] ) );
  INVX1 U14 ( .A(B[28]), .Y(\B_not[28] ) );
  INVX1 U15 ( .A(B[27]), .Y(\B_not[27] ) );
  INVX1 U16 ( .A(B[26]), .Y(\B_not[26] ) );
  INVX1 U17 ( .A(B[25]), .Y(\B_not[25] ) );
  INVX1 U18 ( .A(B[24]), .Y(\B_not[24] ) );
  INVX1 U19 ( .A(B[23]), .Y(\B_not[23] ) );
  INVX1 U20 ( .A(B[22]), .Y(\B_not[22] ) );
  INVX1 U21 ( .A(B[21]), .Y(\B_not[21] ) );
  INVX1 U22 ( .A(B[20]), .Y(\B_not[20] ) );
  INVX1 U23 ( .A(B[1]), .Y(\B_not[1] ) );
  INVX1 U24 ( .A(B[19]), .Y(\B_not[19] ) );
  INVX1 U25 ( .A(B[18]), .Y(\B_not[18] ) );
  INVX1 U26 ( .A(B[17]), .Y(\B_not[17] ) );
  INVX1 U27 ( .A(B[16]), .Y(\B_not[16] ) );
  INVX1 U28 ( .A(B[15]), .Y(\B_not[15] ) );
  INVX1 U29 ( .A(B[14]), .Y(\B_not[14] ) );
  INVX1 U30 ( .A(B[13]), .Y(\B_not[13] ) );
  INVX1 U31 ( .A(B[12]), .Y(\B_not[12] ) );
  INVX1 U32 ( .A(B[11]), .Y(\B_not[11] ) );
  INVX1 U33 ( .A(B[10]), .Y(\B_not[10] ) );
  INVX1 U34 ( .A(B[0]), .Y(\B_not[0] ) );
endmodule


module ALU_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188;

  NAND2X1 U3 ( .A(n188), .B(SH[1]), .Y(n1) );
  NAND2X1 U4 ( .A(SH[0]), .B(SH[1]), .Y(n2) );
  INVX1 U5 ( .A(n135), .Y(n81) );
  INVX1 U6 ( .A(n140), .Y(n12) );
  NAND2X1 U7 ( .A(n81), .B(n159), .Y(n6) );
  INVX1 U8 ( .A(n159), .Y(n77) );
  INVX1 U9 ( .A(n59), .Y(n3) );
  INVX1 U10 ( .A(n60), .Y(n4) );
  NOR2X1 U11 ( .A(n184), .B(SH[3]), .Y(n53) );
  NOR2BX1 U12 ( .AN(n157), .B(SH[2]), .Y(n14) );
  NOR2X1 U13 ( .A(SH[2]), .B(n161), .Y(n55) );
  NAND2BX1 U14 ( .AN(n47), .B(SH[4]), .Y(n8) );
  OAI221XL U15 ( .A0(n5), .A1(n6), .B0(n7), .B1(n8), .C0(n9), .Y(B[9]) );
  AOI222X1 U16 ( .A0(n10), .A1(n11), .B0(n12), .B1(n13), .C0(n14), .C1(n15), 
        .Y(n9) );
  INVX1 U17 ( .A(n16), .Y(n5) );
  OAI221XL U18 ( .A0(n17), .A1(n6), .B0(n18), .B1(n8), .C0(n19), .Y(B[8]) );
  AOI222X1 U19 ( .A0(n10), .A1(n20), .B0(n12), .B1(n21), .C0(n14), .C1(n22), 
        .Y(n19) );
  INVX1 U20 ( .A(n23), .Y(n17) );
  OAI221XL U21 ( .A0(n24), .A1(n6), .B0(n25), .B1(n8), .C0(n26), .Y(B[7]) );
  AOI222X1 U22 ( .A0(n10), .A1(n27), .B0(n12), .B1(n28), .C0(n14), .C1(n29), 
        .Y(n26) );
  INVX1 U23 ( .A(n30), .Y(n24) );
  OAI221XL U24 ( .A0(n31), .A1(n6), .B0(n32), .B1(n8), .C0(n33), .Y(B[6]) );
  AOI222X1 U25 ( .A0(n10), .A1(n34), .B0(n12), .B1(n35), .C0(n14), .C1(n36), 
        .Y(n33) );
  INVX1 U26 ( .A(n37), .Y(n31) );
  OAI221XL U27 ( .A0(n38), .A1(n6), .B0(n39), .B1(n8), .C0(n40), .Y(B[5]) );
  AOI222X1 U28 ( .A0(n10), .A1(n15), .B0(n12), .B1(n16), .C0(n14), .C1(n13), 
        .Y(n40) );
  INVX1 U29 ( .A(n41), .Y(n38) );
  OAI221XL U30 ( .A0(n42), .A1(n6), .B0(n43), .B1(n8), .C0(n44), .Y(B[4]) );
  AOI222X1 U31 ( .A0(n10), .A1(n22), .B0(n12), .B1(n23), .C0(n14), .C1(n21), 
        .Y(n44) );
  INVX1 U32 ( .A(n45), .Y(n42) );
  NOR2X1 U33 ( .A(n46), .B(n47), .Y(B[3]) );
  AOI21X1 U34 ( .A0(n48), .A1(n49), .B0(n50), .Y(n46) );
  MXI2X1 U35 ( .A(n51), .B(n52), .S0(SH[4]), .Y(n50) );
  AOI222X1 U36 ( .A0(n53), .A1(n30), .B0(n54), .B1(n29), .C0(n55), .C1(n28), 
        .Y(n51) );
  OAI221XL U37 ( .A0(n2), .A1(n56), .B0(n1), .B1(n57), .C0(n58), .Y(n30) );
  AOI22X1 U38 ( .A0(A[8]), .A1(n59), .B0(A[7]), .B1(n60), .Y(n58) );
  OAI221XL U39 ( .A0(n2), .A1(n61), .B0(n1), .B1(n62), .C0(n63), .Y(n49) );
  AOI22X1 U40 ( .A0(A[4]), .A1(n59), .B0(A[3]), .B1(n60), .Y(n63) );
  NOR2BX1 U41 ( .AN(n64), .B(n6), .Y(B[31]) );
  NOR2X1 U42 ( .A(n65), .B(n6), .Y(B[30]) );
  NOR2X1 U43 ( .A(n66), .B(n47), .Y(B[2]) );
  AOI21X1 U44 ( .A0(n48), .A1(n67), .B0(n68), .Y(n66) );
  MXI2X1 U45 ( .A(n69), .B(n70), .S0(SH[4]), .Y(n68) );
  AOI222X1 U46 ( .A0(n53), .A1(n37), .B0(n54), .B1(n36), .C0(n55), .C1(n35), 
        .Y(n69) );
  OAI221XL U47 ( .A0(n2), .A1(n57), .B0(n1), .B1(n71), .C0(n72), .Y(n37) );
  AOI22X1 U48 ( .A0(A[7]), .A1(n59), .B0(A[6]), .B1(n60), .Y(n72) );
  INVX1 U49 ( .A(A[9]), .Y(n57) );
  OAI221XL U50 ( .A0(n2), .A1(n62), .B0(n1), .B1(n73), .C0(n74), .Y(n67) );
  AOI22X1 U51 ( .A0(A[3]), .A1(n59), .B0(A[2]), .B1(n60), .Y(n74) );
  INVX1 U52 ( .A(A[5]), .Y(n62) );
  NOR2BX1 U53 ( .AN(n75), .B(n6), .Y(B[29]) );
  NOR2BX1 U54 ( .AN(n76), .B(n6), .Y(B[28]) );
  NOR3X1 U55 ( .A(n77), .B(SH[3]), .C(n78), .Y(B[27]) );
  NOR2X1 U56 ( .A(n79), .B(n77), .Y(B[26]) );
  NOR2X1 U57 ( .A(n7), .B(n77), .Y(B[25]) );
  AOI22X1 U58 ( .A0(n80), .A1(n81), .B0(n75), .B1(n53), .Y(n7) );
  NOR2X1 U59 ( .A(n18), .B(n77), .Y(B[24]) );
  AOI22X1 U60 ( .A0(n82), .A1(n81), .B0(n76), .B1(n53), .Y(n18) );
  NOR2X1 U61 ( .A(n25), .B(n77), .Y(B[23]) );
  AOI222X1 U62 ( .A0(n83), .A1(n53), .B0(n64), .B1(n55), .C0(n84), .C1(n81), 
        .Y(n25) );
  NOR2X1 U63 ( .A(n32), .B(n77), .Y(B[22]) );
  AOI222X1 U64 ( .A0(n85), .A1(n53), .B0(n86), .B1(n55), .C0(n87), .C1(n81), 
        .Y(n32) );
  NOR2X1 U65 ( .A(n39), .B(n77), .Y(B[21]) );
  AOI222X1 U66 ( .A0(n80), .A1(n53), .B0(n75), .B1(n55), .C0(n11), .C1(n81), 
        .Y(n39) );
  NOR2X1 U67 ( .A(n43), .B(n77), .Y(B[20]) );
  AOI222X1 U68 ( .A0(n82), .A1(n53), .B0(n76), .B1(n55), .C0(n20), .C1(n81), 
        .Y(n43) );
  NOR2X1 U69 ( .A(n88), .B(n47), .Y(B[1]) );
  AOI21X1 U70 ( .A0(n48), .A1(n89), .B0(n90), .Y(n88) );
  MXI2X1 U71 ( .A(n91), .B(n92), .S0(SH[4]), .Y(n90) );
  AOI222X1 U72 ( .A0(n53), .A1(n41), .B0(n54), .B1(n13), .C0(n55), .C1(n16), 
        .Y(n91) );
  OAI221XL U73 ( .A0(n2), .A1(n93), .B0(n1), .B1(n94), .C0(n95), .Y(n16) );
  AOI22X1 U74 ( .A0(A[10]), .A1(n59), .B0(A[9]), .B1(n60), .Y(n95) );
  OAI221XL U75 ( .A0(n2), .A1(n71), .B0(n1), .B1(n96), .C0(n97), .Y(n41) );
  AOI22X1 U76 ( .A0(A[6]), .A1(n59), .B0(A[5]), .B1(n60), .Y(n97) );
  INVX1 U77 ( .A(A[8]), .Y(n71) );
  OAI221XL U78 ( .A0(n2), .A1(n73), .B0(n1), .B1(n98), .C0(n99), .Y(n89) );
  AOI22X1 U79 ( .A0(A[2]), .A1(n59), .B0(A[1]), .B1(n60), .Y(n99) );
  INVX1 U80 ( .A(A[4]), .Y(n73) );
  NOR2X1 U81 ( .A(n52), .B(n77), .Y(B[19]) );
  AOI222X1 U82 ( .A0(n27), .A1(n81), .B0(n84), .B1(n53), .C0(SH[3]), .C1(n100), 
        .Y(n52) );
  INVX1 U83 ( .A(n78), .Y(n100) );
  NOR2X1 U84 ( .A(n70), .B(n77), .Y(B[18]) );
  AOI221X1 U85 ( .A0(n87), .A1(n53), .B0(n34), .B1(n81), .C0(n101), .Y(n70) );
  INVX1 U86 ( .A(n102), .Y(n101) );
  AOI22X1 U87 ( .A0(n54), .A1(n86), .B0(n55), .B1(n85), .Y(n102) );
  NOR2X1 U88 ( .A(n92), .B(n77), .Y(B[17]) );
  AOI221X1 U89 ( .A0(n11), .A1(n53), .B0(n15), .B1(n81), .C0(n103), .Y(n92) );
  INVX1 U90 ( .A(n104), .Y(n103) );
  AOI22X1 U91 ( .A0(n54), .A1(n75), .B0(n55), .B1(n80), .Y(n104) );
  NOR2X1 U92 ( .A(n105), .B(n77), .Y(B[16]) );
  OAI221XL U93 ( .A0(n106), .A1(n107), .B0(n108), .B1(n6), .C0(n109), .Y(B[15]) );
  AOI222X1 U94 ( .A0(n14), .A1(n84), .B0(n110), .B1(n64), .C0(n12), .C1(n27), 
        .Y(n109) );
  INVX1 U95 ( .A(n83), .Y(n106) );
  OAI221XL U96 ( .A0(n111), .A1(n107), .B0(n112), .B1(n6), .C0(n113), .Y(B[14]) );
  AOI222X1 U97 ( .A0(n14), .A1(n87), .B0(n110), .B1(n86), .C0(n12), .C1(n34), 
        .Y(n113) );
  INVX1 U98 ( .A(n36), .Y(n112) );
  INVX1 U99 ( .A(n85), .Y(n111) );
  OAI221XL U100 ( .A0(n114), .A1(n107), .B0(n115), .B1(n6), .C0(n116), .Y(
        B[13]) );
  AOI222X1 U101 ( .A0(n14), .A1(n11), .B0(n110), .B1(n75), .C0(n12), .C1(n15), 
        .Y(n116) );
  OAI221XL U102 ( .A0(n2), .A1(n117), .B0(n1), .B1(n118), .C0(n119), .Y(n15)
         );
  AOI22X1 U103 ( .A0(A[18]), .A1(n59), .B0(A[17]), .B1(n60), .Y(n119) );
  OAI222XL U104 ( .A0(n3), .A1(n120), .B0(n1), .B1(n121), .C0(n4), .C1(n122), 
        .Y(n75) );
  OAI221XL U105 ( .A0(n2), .A1(n123), .B0(n1), .B1(n124), .C0(n125), .Y(n11)
         );
  AOI22X1 U106 ( .A0(A[22]), .A1(n59), .B0(A[21]), .B1(n60), .Y(n125) );
  INVX1 U107 ( .A(n13), .Y(n115) );
  OAI221XL U108 ( .A0(n2), .A1(n126), .B0(n1), .B1(n127), .C0(n128), .Y(n13)
         );
  AOI22X1 U109 ( .A0(A[14]), .A1(n59), .B0(A[13]), .B1(n60), .Y(n128) );
  INVX1 U110 ( .A(n80), .Y(n114) );
  OAI221XL U111 ( .A0(n2), .A1(n129), .B0(n1), .B1(n130), .C0(n131), .Y(n80)
         );
  AOI22X1 U112 ( .A0(A[26]), .A1(n59), .B0(A[25]), .B1(n60), .Y(n131) );
  OAI221XL U113 ( .A0(n132), .A1(n107), .B0(n133), .B1(n6), .C0(n134), .Y(
        B[12]) );
  AOI222X1 U114 ( .A0(n14), .A1(n20), .B0(n110), .B1(n76), .C0(n12), .C1(n22), 
        .Y(n134) );
  NOR2X1 U115 ( .A(n8), .B(n135), .Y(n110) );
  INVX1 U116 ( .A(n21), .Y(n133) );
  INVX1 U117 ( .A(n82), .Y(n132) );
  OAI221XL U118 ( .A0(n136), .A1(n107), .B0(n137), .B1(n6), .C0(n138), .Y(
        B[11]) );
  AOI21X1 U119 ( .A0(n14), .A1(n27), .B0(n139), .Y(n138) );
  OAI32X1 U120 ( .A0(n8), .A1(SH[3]), .A2(n78), .B0(n108), .B1(n140), .Y(n139)
         );
  INVX1 U121 ( .A(n29), .Y(n108) );
  OAI221XL U122 ( .A0(n2), .A1(n141), .B0(n1), .B1(n142), .C0(n143), .Y(n29)
         );
  AOI22X1 U123 ( .A0(n59), .A1(A[16]), .B0(n60), .B1(A[15]), .Y(n143) );
  MXI2X1 U124 ( .A(n83), .B(n64), .S0(SH[2]), .Y(n78) );
  NOR2X1 U125 ( .A(n121), .B(n4), .Y(n64) );
  OAI221XL U126 ( .A0(n2), .A1(n120), .B0(n1), .B1(n122), .C0(n144), .Y(n83)
         );
  AOI22X1 U127 ( .A0(A[28]), .A1(n59), .B0(A[27]), .B1(n60), .Y(n144) );
  OAI221XL U128 ( .A0(n2), .A1(n145), .B0(n1), .B1(n146), .C0(n147), .Y(n27)
         );
  AOI22X1 U129 ( .A0(A[20]), .A1(n59), .B0(A[19]), .B1(n60), .Y(n147) );
  INVX1 U130 ( .A(n28), .Y(n137) );
  OAI221XL U131 ( .A0(n2), .A1(n148), .B0(n1), .B1(n149), .C0(n150), .Y(n28)
         );
  AOI22X1 U132 ( .A0(A[12]), .A1(n59), .B0(A[11]), .B1(n60), .Y(n150) );
  INVX1 U133 ( .A(n84), .Y(n136) );
  OAI221XL U134 ( .A0(n2), .A1(n151), .B0(n1), .B1(n152), .C0(n153), .Y(n84)
         );
  AOI22X1 U135 ( .A0(A[24]), .A1(n59), .B0(A[23]), .B1(n60), .Y(n153) );
  OAI221XL U136 ( .A0(n154), .A1(n6), .B0(n79), .B1(n8), .C0(n155), .Y(B[10])
         );
  AOI222X1 U137 ( .A0(n10), .A1(n87), .B0(n12), .B1(n36), .C0(n14), .C1(n34), 
        .Y(n155) );
  OAI221XL U138 ( .A0(n2), .A1(n146), .B0(n1), .B1(n117), .C0(n156), .Y(n34)
         );
  AOI22X1 U139 ( .A0(A[19]), .A1(n59), .B0(A[18]), .B1(n60), .Y(n156) );
  INVX1 U140 ( .A(A[20]), .Y(n117) );
  INVX1 U141 ( .A(A[21]), .Y(n146) );
  OAI221XL U142 ( .A0(n2), .A1(n142), .B0(n126), .B1(n1), .C0(n158), .Y(n36)
         );
  AOI22X1 U143 ( .A0(n59), .A1(A[15]), .B0(n60), .B1(A[14]), .Y(n158) );
  INVX1 U144 ( .A(A[16]), .Y(n126) );
  INVX1 U145 ( .A(A[17]), .Y(n142) );
  NAND2X1 U146 ( .A(n159), .B(n53), .Y(n140) );
  OAI221XL U147 ( .A0(n2), .A1(n152), .B0(n1), .B1(n123), .C0(n160), .Y(n87)
         );
  AOI22X1 U148 ( .A0(A[23]), .A1(n59), .B0(A[22]), .B1(n60), .Y(n160) );
  INVX1 U149 ( .A(A[24]), .Y(n123) );
  INVX1 U150 ( .A(A[25]), .Y(n152) );
  INVX1 U151 ( .A(n107), .Y(n10) );
  NAND2X1 U152 ( .A(n157), .B(SH[2]), .Y(n107) );
  NOR2X1 U153 ( .A(n77), .B(n161), .Y(n157) );
  AOI22X1 U154 ( .A0(n85), .A1(n81), .B0(n86), .B1(n53), .Y(n79) );
  INVX1 U155 ( .A(n65), .Y(n86) );
  AOI22X1 U156 ( .A0(n60), .A1(A[30]), .B0(n59), .B1(A[31]), .Y(n65) );
  OAI221XL U157 ( .A0(n2), .A1(n122), .B0(n1), .B1(n129), .C0(n162), .Y(n85)
         );
  AOI22X1 U158 ( .A0(A[27]), .A1(n59), .B0(A[26]), .B1(n60), .Y(n162) );
  INVX1 U159 ( .A(A[28]), .Y(n129) );
  INVX1 U160 ( .A(A[29]), .Y(n122) );
  NOR2X1 U161 ( .A(n47), .B(SH[4]), .Y(n159) );
  INVX1 U162 ( .A(n35), .Y(n154) );
  OAI221XL U163 ( .A0(n2), .A1(n149), .B0(n1), .B1(n93), .C0(n163), .Y(n35) );
  AOI22X1 U164 ( .A0(A[11]), .A1(n59), .B0(A[10]), .B1(n60), .Y(n163) );
  INVX1 U165 ( .A(A[12]), .Y(n93) );
  INVX1 U166 ( .A(A[13]), .Y(n149) );
  NOR2X1 U167 ( .A(n164), .B(n47), .Y(B[0]) );
  NAND4X1 U168 ( .A(n165), .B(n166), .C(n167), .D(n168), .Y(n47) );
  NOR4BX1 U169 ( .AN(n169), .B(SH[5]), .C(SH[30]), .D(SH[31]), .Y(n168) );
  NOR4X1 U170 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n169) );
  NOR4BX1 U171 ( .AN(n170), .B(SH[25]), .C(SH[23]), .D(SH[24]), .Y(n167) );
  NOR4X1 U172 ( .A(SH[29]), .B(SH[28]), .C(SH[27]), .D(SH[26]), .Y(n170) );
  NOR4BX1 U173 ( .AN(n171), .B(SH[18]), .C(SH[16]), .D(SH[17]), .Y(n166) );
  NOR4X1 U174 ( .A(SH[22]), .B(SH[21]), .C(SH[20]), .D(SH[19]), .Y(n171) );
  NOR4BX1 U175 ( .AN(n172), .B(SH[12]), .C(SH[10]), .D(SH[11]), .Y(n165) );
  NOR3X1 U176 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n172) );
  AOI21X1 U177 ( .A0(n48), .A1(n173), .B0(n174), .Y(n164) );
  MXI2X1 U178 ( .A(n175), .B(n105), .S0(SH[4]), .Y(n174) );
  AOI221X1 U179 ( .A0(n20), .A1(n53), .B0(n22), .B1(n81), .C0(n176), .Y(n105)
         );
  INVX1 U180 ( .A(n177), .Y(n176) );
  AOI22X1 U181 ( .A0(n54), .A1(n76), .B0(n55), .B1(n82), .Y(n177) );
  OAI221XL U182 ( .A0(n2), .A1(n130), .B0(n1), .B1(n151), .C0(n178), .Y(n82)
         );
  AOI22X1 U183 ( .A0(A[25]), .A1(n59), .B0(A[24]), .B1(n60), .Y(n178) );
  INVX1 U184 ( .A(A[26]), .Y(n151) );
  INVX1 U185 ( .A(A[27]), .Y(n130) );
  OAI221XL U186 ( .A0(n2), .A1(n121), .B0(n1), .B1(n120), .C0(n179), .Y(n76)
         );
  AOI22X1 U187 ( .A0(A[29]), .A1(n59), .B0(A[28]), .B1(n60), .Y(n179) );
  INVX1 U188 ( .A(A[30]), .Y(n120) );
  INVX1 U189 ( .A(A[31]), .Y(n121) );
  OAI221XL U190 ( .A0(n2), .A1(n118), .B0(n1), .B1(n141), .C0(n180), .Y(n22)
         );
  AOI22X1 U191 ( .A0(A[17]), .A1(n59), .B0(n60), .B1(A[16]), .Y(n180) );
  INVX1 U192 ( .A(A[18]), .Y(n141) );
  INVX1 U193 ( .A(A[19]), .Y(n118) );
  OAI221XL U194 ( .A0(n2), .A1(n124), .B0(n1), .B1(n145), .C0(n181), .Y(n20)
         );
  AOI22X1 U195 ( .A0(A[21]), .A1(n59), .B0(A[20]), .B1(n60), .Y(n181) );
  INVX1 U196 ( .A(A[22]), .Y(n145) );
  INVX1 U197 ( .A(A[23]), .Y(n124) );
  AOI222X1 U198 ( .A0(n53), .A1(n45), .B0(n54), .B1(n21), .C0(n55), .C1(n23), 
        .Y(n175) );
  OAI221XL U199 ( .A0(n2), .A1(n94), .B0(n1), .B1(n56), .C0(n182), .Y(n23) );
  AOI22X1 U200 ( .A0(A[9]), .A1(n59), .B0(A[8]), .B1(n60), .Y(n182) );
  INVX1 U201 ( .A(A[10]), .Y(n56) );
  INVX1 U202 ( .A(A[11]), .Y(n94) );
  OAI221XL U203 ( .A0(n2), .A1(n127), .B0(n1), .B1(n148), .C0(n183), .Y(n21)
         );
  AOI22X1 U204 ( .A0(A[13]), .A1(n59), .B0(A[12]), .B1(n60), .Y(n183) );
  INVX1 U205 ( .A(A[14]), .Y(n148) );
  INVX1 U206 ( .A(A[15]), .Y(n127) );
  NOR2X1 U207 ( .A(n184), .B(n161), .Y(n54) );
  OAI221XL U208 ( .A0(n2), .A1(n96), .B0(n1), .B1(n61), .C0(n185), .Y(n45) );
  AOI22X1 U209 ( .A0(A[5]), .A1(n59), .B0(A[4]), .B1(n60), .Y(n185) );
  INVX1 U210 ( .A(A[6]), .Y(n61) );
  INVX1 U211 ( .A(A[7]), .Y(n96) );
  OAI221XL U212 ( .A0(n2), .A1(n98), .B0(n1), .B1(n186), .C0(n187), .Y(n173)
         );
  AOI22X1 U213 ( .A0(A[1]), .A1(n59), .B0(A[0]), .B1(n60), .Y(n187) );
  NOR2X1 U214 ( .A(SH[0]), .B(SH[1]), .Y(n60) );
  NOR2X1 U215 ( .A(n188), .B(SH[1]), .Y(n59) );
  INVX1 U216 ( .A(A[2]), .Y(n186) );
  INVX1 U217 ( .A(SH[0]), .Y(n188) );
  INVX1 U218 ( .A(A[3]), .Y(n98) );
  NOR2X1 U219 ( .A(n135), .B(SH[4]), .Y(n48) );
  NAND2X1 U220 ( .A(n184), .B(n161), .Y(n135) );
  INVX1 U221 ( .A(SH[3]), .Y(n161) );
  INVX1 U222 ( .A(SH[2]), .Y(n184) );
endmodule


module ALU_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \SHMAG[5] , \SHMAG[4] , \SHMAG[3] , \SHMAG[2] , \SHMAG[1] ,
         \SHMAG[0] , \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] ,
         \ML_int[1][28] , \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] ,
         \ML_int[1][24] , \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] ,
         \ML_int[1][20] , \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] ,
         \ML_int[1][16] , \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] ,
         \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] ,
         \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] ,
         \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] ,
         \ML_int[1][0] , \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] ,
         \ML_int[2][28] , \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] ,
         \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] ,
         \ML_int[2][20] , \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] ,
         \ML_int[2][16] , \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] ,
         \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] ,
         \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] ,
         \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] ,
         \ML_int[2][0] , \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] ,
         \ML_int[3][28] , \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] ,
         \ML_int[3][24] , \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] ,
         \ML_int[3][20] , \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] ,
         \ML_int[3][16] , \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] ,
         \ML_int[3][12] , \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] ,
         \ML_int[3][8] , \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] ,
         \ML_int[3][4] , \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] ,
         \ML_int[3][0] , \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] ,
         \ML_int[4][28] , \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] ,
         \ML_int[4][24] , \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] ,
         \ML_int[4][20] , \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] ,
         \ML_int[4][16] , \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] ,
         \ML_int[4][12] , \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] ,
         \ML_int[4][4] , \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] ,
         \ML_int[4][0] , \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] ,
         \ML_int[5][28] , \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] ,
         \ML_int[5][24] , \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] ,
         \ML_int[5][20] , \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] ,
         \ML_int[5][16] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38;

  MX2X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S0(n1), .Y(\ML_int[1][31] ) );
  MX2X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S0(n2), .Y(
        \ML_int[2][31] ) );
  MX2X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S0(n3), .Y(
        \ML_int[3][31] ) );
  MX2X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S0(n4), .Y(
        \ML_int[4][31] ) );
  MX2X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S0(n1), .Y(\ML_int[1][30] ) );
  MX2X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S0(n2), .Y(
        \ML_int[2][30] ) );
  MX2X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S0(n3), .Y(
        \ML_int[3][30] ) );
  MX2X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S0(n1), .Y(\ML_int[1][1] ) );
  MX2X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S0(n1), .Y(\ML_int[1][2] ) );
  MX2X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S0(n1), .Y(\ML_int[1][27] ) );
  MX2X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S0(n1), .Y(\ML_int[1][25] ) );
  MX2X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S0(n1), .Y(\ML_int[1][29] ) );
  MX2X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S0(n1), .Y(\ML_int[1][23] ) );
  MX2X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S0(n1), .Y(\ML_int[1][21] ) );
  MX2X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S0(n1), .Y(\ML_int[1][19] ) );
  MX2X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S0(n1), .Y(\ML_int[1][17] ) );
  MX2X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S0(n1), .Y(\ML_int[1][26] ) );
  MX2X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S0(n1), .Y(\ML_int[1][24] ) );
  MX2X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S0(n1), .Y(\ML_int[1][28] ) );
  MX2X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S0(n1), .Y(\ML_int[1][22] ) );
  MX2X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S0(n1), .Y(\ML_int[1][20] ) );
  MX2X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S0(n1), .Y(\ML_int[1][18] ) );
  MX2X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S0(n1), .Y(\ML_int[1][16] ) );
  MX2X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S0(n1), .Y(\ML_int[1][15] ) );
  MX2X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S0(n1), .Y(\ML_int[1][14] ) );
  MX2X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S0(n1), .Y(\ML_int[1][13] ) );
  MX2X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S0(n1), .Y(\ML_int[1][12] ) );
  MX2X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S0(n1), .Y(\ML_int[1][11] ) );
  MX2X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S0(n1), .Y(\ML_int[1][10] ) );
  MX2X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S0(n1), .Y(\ML_int[1][9] ) );
  MX2X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S0(n1), .Y(\ML_int[1][8] ) );
  MX2X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S0(n1), .Y(\ML_int[1][7] ) );
  MX2X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S0(n1), .Y(\ML_int[1][5] ) );
  MX2X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S0(n1), .Y(\ML_int[1][3] ) );
  MX2X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S0(n1), .Y(\ML_int[1][6] ) );
  MX2X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S0(n1), .Y(\ML_int[1][4] ) );
  MX2X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S0(n5), .Y(
        \ML_int[5][31] ) );
  MX2X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S0(n2), .Y(
        \ML_int[2][29] ) );
  MX2X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S0(n3), .Y(
        \ML_int[3][29] ) );
  MX2X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S0(n2), .Y(
        \ML_int[2][28] ) );
  MX2X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S0(n3), .Y(
        \ML_int[3][28] ) );
  MX2X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S0(n2), .Y(
        \ML_int[2][3] ) );
  MX2X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S0(n2), .Y(
        \ML_int[2][2] ) );
  MX2X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S0(n2), .Y(
        \ML_int[2][9] ) );
  MX2X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S0(n2), .Y(
        \ML_int[2][27] ) );
  MX2X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S0(n2), .Y(
        \ML_int[2][23] ) );
  MX2X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S0(n2), .Y(
        \ML_int[2][19] ) );
  MX2X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S0(n2), .Y(
        \ML_int[2][26] ) );
  MX2X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S0(n2), .Y(
        \ML_int[2][22] ) );
  MX2X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S0(n2), .Y(
        \ML_int[2][18] ) );
  MX2X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S0(n2), .Y(
        \ML_int[2][25] ) );
  MX2X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S0(n2), .Y(
        \ML_int[2][21] ) );
  MX2X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S0(n2), .Y(
        \ML_int[2][17] ) );
  MX2X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S0(n2), .Y(
        \ML_int[2][24] ) );
  MX2X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S0(n2), .Y(
        \ML_int[2][16] ) );
  MX2X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S0(n2), .Y(
        \ML_int[2][20] ) );
  MX2X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S0(n2), .Y(
        \ML_int[2][15] ) );
  MX2X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S0(n2), .Y(
        \ML_int[2][14] ) );
  MX2X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S0(n2), .Y(
        \ML_int[2][13] ) );
  MX2X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S0(n2), .Y(
        \ML_int[2][12] ) );
  MX2X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S0(n2), .Y(
        \ML_int[2][11] ) );
  MX2X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S0(n2), .Y(
        \ML_int[2][10] ) );
  MX2X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S0(n2), .Y(
        \ML_int[2][8] ) );
  MX2X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S0(n2), .Y(
        \ML_int[2][7] ) );
  MX2X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S0(n2), .Y(
        \ML_int[2][6] ) );
  MX2X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S0(n2), .Y(
        \ML_int[2][5] ) );
  MX2X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S0(n2), .Y(
        \ML_int[2][4] ) );
  MX2X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S0(n4), .Y(
        \ML_int[4][16] ) );
  MX2X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S0(n5), .Y(
        \ML_int[5][16] ) );
  MX2X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S0(n5), .Y(
        \ML_int[5][20] ) );
  MX2X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S0(n4), .Y(
        \ML_int[4][19] ) );
  MX2X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S0(n5), .Y(
        \ML_int[5][19] ) );
  MX2X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S0(n4), .Y(
        \ML_int[4][18] ) );
  MX2X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S0(n5), .Y(
        \ML_int[5][18] ) );
  MX2X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S0(n4), .Y(
        \ML_int[4][17] ) );
  MX2X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S0(n5), .Y(
        \ML_int[5][17] ) );
  MX2X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S0(n4), .Y(
        \ML_int[4][30] ) );
  MX2X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S0(n5), .Y(
        \ML_int[5][30] ) );
  MX2X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S0(n4), .Y(
        \ML_int[4][29] ) );
  MX2X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S0(n5), .Y(
        \ML_int[5][29] ) );
  MX2X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S0(n4), .Y(
        \ML_int[4][28] ) );
  MX2X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S0(n5), .Y(
        \ML_int[5][28] ) );
  MX2X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S0(n4), .Y(
        \ML_int[4][27] ) );
  MX2X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S0(n5), .Y(
        \ML_int[5][27] ) );
  MX2X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S0(n4), .Y(
        \ML_int[4][26] ) );
  MX2X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S0(n5), .Y(
        \ML_int[5][26] ) );
  MX2X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S0(n4), .Y(
        \ML_int[4][25] ) );
  MX2X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S0(n5), .Y(
        \ML_int[5][25] ) );
  MX2X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S0(n4), .Y(
        \ML_int[4][24] ) );
  MX2X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S0(n5), .Y(
        \ML_int[5][24] ) );
  MX2X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S0(n5), .Y(
        \ML_int[5][23] ) );
  MX2X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S0(n5), .Y(
        \ML_int[5][22] ) );
  MX2X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S0(n4), .Y(
        \ML_int[4][21] ) );
  MX2X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S0(n5), .Y(
        \ML_int[5][21] ) );
  MX2X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S0(n3), .Y(
        \ML_int[3][27] ) );
  MX2X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S0(n3), .Y(
        \ML_int[3][26] ) );
  MX2X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S0(n3), .Y(
        \ML_int[3][25] ) );
  MX2X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S0(n3), .Y(
        \ML_int[3][24] ) );
  MX2X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S0(n3), .Y(
        \ML_int[3][7] ) );
  MX2X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S0(n3), .Y(
        \ML_int[3][6] ) );
  MX2X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S0(n3), .Y(
        \ML_int[3][5] ) );
  MX2X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S0(n3), .Y(
        \ML_int[3][4] ) );
  MX2X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S0(n3), .Y(
        \ML_int[3][13] ) );
  MX2X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S0(n3), .Y(
        \ML_int[3][11] ) );
  MX2X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S0(n3), .Y(
        \ML_int[3][10] ) );
  MX2X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S0(n3), .Y(
        \ML_int[3][9] ) );
  MX2X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S0(n3), .Y(
        \ML_int[3][8] ) );
  MX2X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S0(n3), .Y(
        \ML_int[3][23] ) );
  MX2X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S0(n3), .Y(
        \ML_int[3][21] ) );
  MX2X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S0(n3), .Y(
        \ML_int[3][20] ) );
  MX2X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S0(n3), .Y(
        \ML_int[3][19] ) );
  MX2X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S0(n3), .Y(
        \ML_int[3][18] ) );
  MX2X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S0(n3), .Y(
        \ML_int[3][17] ) );
  MX2X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S0(n3), .Y(
        \ML_int[3][16] ) );
  MX2X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S0(n3), .Y(
        \ML_int[3][15] ) );
  MX2X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S0(n3), .Y(
        \ML_int[3][14] ) );
  MX2X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S0(n3), .Y(
        \ML_int[3][12] ) );
  MX2X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S0(n4), .Y(
        \ML_int[4][23] ) );
  MX2X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S0(n4), .Y(
        \ML_int[4][22] ) );
  MX2X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S0(n4), .Y(
        \ML_int[4][20] ) );
  MX2X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S0(n4), .Y(
        \ML_int[4][15] ) );
  MX2X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S0(n4), .Y(
        \ML_int[4][14] ) );
  MX2X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S0(n4), .Y(
        \ML_int[4][13] ) );
  MX2X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S0(n4), .Y(
        \ML_int[4][12] ) );
  MX2X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S0(n4), .Y(
        \ML_int[4][11] ) );
  MX2X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S0(n4), .Y(
        \ML_int[4][10] ) );
  MX2X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S0(n4), .Y(
        \ML_int[4][9] ) );
  MX2X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S0(n4), .Y(
        \ML_int[4][8] ) );
  INVX1 U3 ( .A(\SHMAG[1] ), .Y(n2) );
  INVX1 U4 ( .A(\SHMAG[2] ), .Y(n3) );
  INVX1 U5 ( .A(\SHMAG[3] ), .Y(n4) );
  INVX1 U6 ( .A(\SHMAG[4] ), .Y(n5) );
  MX2X1 U7 ( .A(\ML_int[2][18] ), .B(\ML_int[2][22] ), .S0(\SHMAG[2] ), .Y(
        \ML_int[3][22] ) );
  INVX1 U8 ( .A(\SHMAG[0] ), .Y(n1) );
  OR2X2 U9 ( .A(n13), .B(n5), .Y(n7) );
  NAND2BX1 U10 ( .AN(n6), .B(n19), .Y(n13) );
  INVX1 U11 ( .A(\SHMAG[5] ), .Y(n6) );
  NOR2BX1 U12 ( .AN(\ML_int[4][9] ), .B(n7), .Y(B[9]) );
  NOR2BX1 U13 ( .AN(\ML_int[4][8] ), .B(n7), .Y(B[8]) );
  NOR2X1 U14 ( .A(n7), .B(n8), .Y(B[7]) );
  NOR2X1 U15 ( .A(n7), .B(n9), .Y(B[6]) );
  NOR2X1 U16 ( .A(n7), .B(n10), .Y(B[5]) );
  NOR2X1 U17 ( .A(n7), .B(n11), .Y(B[4]) );
  NOR2X1 U18 ( .A(n7), .B(n12), .Y(B[3]) );
  NOR2BX1 U19 ( .AN(\ML_int[5][31] ), .B(n13), .Y(B[31]) );
  NOR2BX1 U20 ( .AN(\ML_int[5][30] ), .B(n13), .Y(B[30]) );
  NOR2X1 U21 ( .A(n7), .B(n14), .Y(B[2]) );
  NOR2BX1 U22 ( .AN(\ML_int[5][29] ), .B(n13), .Y(B[29]) );
  NOR2BX1 U23 ( .AN(\ML_int[5][28] ), .B(n13), .Y(B[28]) );
  NOR2BX1 U24 ( .AN(\ML_int[5][27] ), .B(n13), .Y(B[27]) );
  NOR2BX1 U25 ( .AN(\ML_int[5][26] ), .B(n13), .Y(B[26]) );
  NOR2BX1 U26 ( .AN(\ML_int[5][25] ), .B(n13), .Y(B[25]) );
  NOR2BX1 U27 ( .AN(\ML_int[5][24] ), .B(n13), .Y(B[24]) );
  NOR2BX1 U28 ( .AN(\ML_int[5][23] ), .B(n13), .Y(B[23]) );
  NOR2BX1 U29 ( .AN(\ML_int[5][22] ), .B(n13), .Y(B[22]) );
  NOR2BX1 U30 ( .AN(\ML_int[5][21] ), .B(n13), .Y(B[21]) );
  NOR2BX1 U31 ( .AN(\ML_int[5][20] ), .B(n13), .Y(B[20]) );
  NOR2X1 U32 ( .A(n7), .B(n15), .Y(B[1]) );
  NOR2BX1 U33 ( .AN(\ML_int[5][19] ), .B(n13), .Y(B[19]) );
  NOR2BX1 U34 ( .AN(\ML_int[5][18] ), .B(n13), .Y(B[18]) );
  NOR2BX1 U35 ( .AN(\ML_int[5][17] ), .B(n13), .Y(B[17]) );
  NOR2BX1 U36 ( .AN(\ML_int[5][16] ), .B(n13), .Y(B[16]) );
  NOR2BX1 U37 ( .AN(\ML_int[4][15] ), .B(n7), .Y(B[15]) );
  NOR2BX1 U38 ( .AN(\ML_int[4][14] ), .B(n7), .Y(B[14]) );
  NOR2BX1 U39 ( .AN(\ML_int[4][13] ), .B(n7), .Y(B[13]) );
  NOR2BX1 U40 ( .AN(\ML_int[4][12] ), .B(n7), .Y(B[12]) );
  NOR2BX1 U41 ( .AN(\ML_int[4][11] ), .B(n7), .Y(B[11]) );
  NOR2BX1 U42 ( .AN(\ML_int[4][10] ), .B(n7), .Y(B[10]) );
  NOR2X1 U43 ( .A(n7), .B(n16), .Y(B[0]) );
  AOI21X1 U44 ( .A0(SH[4]), .A1(n17), .B0(n18), .Y(\SHMAG[4] ) );
  AOI21X1 U45 ( .A0(SH[5]), .A1(n17), .B0(n18), .Y(\SHMAG[5] ) );
  INVX1 U46 ( .A(n8), .Y(\ML_int[4][7] ) );
  NAND2X1 U47 ( .A(\ML_int[3][7] ), .B(\SHMAG[3] ), .Y(n8) );
  INVX1 U48 ( .A(n9), .Y(\ML_int[4][6] ) );
  NAND2X1 U49 ( .A(\ML_int[3][6] ), .B(\SHMAG[3] ), .Y(n9) );
  INVX1 U50 ( .A(n10), .Y(\ML_int[4][5] ) );
  NAND2X1 U51 ( .A(\ML_int[3][5] ), .B(\SHMAG[3] ), .Y(n10) );
  INVX1 U52 ( .A(n11), .Y(\ML_int[4][4] ) );
  NAND2X1 U53 ( .A(\ML_int[3][4] ), .B(\SHMAG[3] ), .Y(n11) );
  INVX1 U54 ( .A(n12), .Y(\ML_int[4][3] ) );
  NAND2X1 U55 ( .A(\ML_int[3][3] ), .B(\SHMAG[3] ), .Y(n12) );
  INVX1 U56 ( .A(n14), .Y(\ML_int[4][2] ) );
  NAND2X1 U57 ( .A(\ML_int[3][2] ), .B(\SHMAG[3] ), .Y(n14) );
  INVX1 U58 ( .A(n15), .Y(\ML_int[4][1] ) );
  NAND2X1 U59 ( .A(\ML_int[3][1] ), .B(\SHMAG[3] ), .Y(n15) );
  INVX1 U60 ( .A(n16), .Y(\ML_int[4][0] ) );
  NAND2X1 U61 ( .A(\ML_int[3][0] ), .B(\SHMAG[3] ), .Y(n16) );
  AOI21X1 U62 ( .A0(SH[3]), .A1(n17), .B0(n18), .Y(\SHMAG[3] ) );
  NOR2BX1 U63 ( .AN(\ML_int[2][3] ), .B(n3), .Y(\ML_int[3][3] ) );
  NOR2BX1 U64 ( .AN(\ML_int[2][2] ), .B(n3), .Y(\ML_int[3][2] ) );
  NOR2BX1 U65 ( .AN(\ML_int[2][1] ), .B(n3), .Y(\ML_int[3][1] ) );
  NOR2BX1 U66 ( .AN(\ML_int[2][0] ), .B(n3), .Y(\ML_int[3][0] ) );
  AOI21X1 U67 ( .A0(SH[2]), .A1(n17), .B0(n18), .Y(\SHMAG[2] ) );
  NOR2BX1 U68 ( .AN(\ML_int[1][1] ), .B(n2), .Y(\ML_int[2][1] ) );
  NOR2BX1 U69 ( .AN(\ML_int[1][0] ), .B(n2), .Y(\ML_int[2][0] ) );
  AOI21X1 U70 ( .A0(SH[1]), .A1(n17), .B0(n18), .Y(\SHMAG[1] ) );
  NOR2BX1 U71 ( .AN(A[0]), .B(n1), .Y(\ML_int[1][0] ) );
  AOI21X1 U72 ( .A0(SH[0]), .A1(n17), .B0(n18), .Y(\SHMAG[0] ) );
  INVX1 U73 ( .A(n20), .Y(n18) );
  OAI31X1 U74 ( .A0(n21), .A1(n22), .A2(n23), .B0(n19), .Y(n20) );
  INVX1 U75 ( .A(SH[31]), .Y(n19) );
  OR4X1 U76 ( .A(n24), .B(SH[11]), .C(SH[12]), .D(SH[10]), .Y(n23) );
  OR3XL U77 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n24) );
  OR4X1 U78 ( .A(n25), .B(SH[17]), .C(SH[18]), .D(SH[16]), .Y(n22) );
  OR3XL U79 ( .A(SH[19]), .B(SH[21]), .C(SH[20]), .Y(n25) );
  NAND4X1 U80 ( .A(n26), .B(n27), .C(n28), .D(n29), .Y(n21) );
  NOR4X1 U81 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n29) );
  NOR3X1 U82 ( .A(SH[28]), .B(SH[30]), .C(SH[29]), .Y(n28) );
  NOR3X1 U83 ( .A(SH[25]), .B(SH[27]), .C(SH[26]), .Y(n27) );
  NOR3X1 U84 ( .A(SH[22]), .B(SH[24]), .C(SH[23]), .Y(n26) );
  OAI31X1 U85 ( .A0(n30), .A1(n31), .A2(n32), .B0(SH[31]), .Y(n17) );
  NAND4X1 U86 ( .A(SH[8]), .B(SH[7]), .C(SH[9]), .D(n33), .Y(n32) );
  AND3X1 U87 ( .A(SH[6]), .B(SH[29]), .C(SH[30]), .Y(n33) );
  NAND4X1 U88 ( .A(SH[27]), .B(SH[26]), .C(SH[28]), .D(n34), .Y(n31) );
  AND3X1 U89 ( .A(SH[25]), .B(SH[23]), .C(SH[24]), .Y(n34) );
  NAND4X1 U90 ( .A(n35), .B(n36), .C(n37), .D(n38), .Y(n30) );
  AND4X1 U91 ( .A(SH[13]), .B(SH[12]), .C(SH[11]), .D(SH[10]), .Y(n38) );
  AND3X1 U92 ( .A(SH[16]), .B(SH[14]), .C(SH[15]), .Y(n37) );
  AND3X1 U93 ( .A(SH[19]), .B(SH[17]), .C(SH[18]), .Y(n36) );
  AND3X1 U94 ( .A(SH[22]), .B(SH[20]), .C(SH[21]), .Y(n35) );
endmodule


module ALU_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] ;

  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        SUM[8]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        SUM[7]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        SUM[6]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        SUM[5]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(\carry[31] ), .Y(SUM[31]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(\carry[1] ) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module CPU_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NOR4BX1 U1 ( .AN(n1), .B(n2), .C(n3), .D(n4), .Y(EQ) );
  NAND4X1 U2 ( .A(n5), .B(n6), .C(n7), .D(n8), .Y(n4) );
  XNOR2X1 U3 ( .A(B[3]), .B(A[3]), .Y(n8) );
  XNOR2X1 U4 ( .A(B[5]), .B(A[5]), .Y(n7) );
  XNOR2X1 U5 ( .A(B[6]), .B(A[6]), .Y(n6) );
  XNOR2X1 U6 ( .A(B[7]), .B(A[7]), .Y(n5) );
  NAND4X1 U7 ( .A(n9), .B(n10), .C(n11), .D(n12), .Y(n3) );
  OAI22X1 U8 ( .A0(n13), .A1(n14), .B0(B[1]), .B1(n13), .Y(n12) );
  INVX1 U9 ( .A(A[1]), .Y(n14) );
  NOR2BX1 U10 ( .AN(B[0]), .B(A[0]), .Y(n13) );
  OAI22X1 U11 ( .A0(A[1]), .A1(n15), .B0(n15), .B1(n16), .Y(n11) );
  INVX1 U12 ( .A(B[1]), .Y(n16) );
  NOR2BX1 U13 ( .AN(A[0]), .B(B[0]), .Y(n15) );
  XNOR2X1 U14 ( .A(B[2]), .B(A[2]), .Y(n10) );
  XNOR2X1 U15 ( .A(B[4]), .B(A[4]), .Y(n9) );
  OR4X1 U16 ( .A(n17), .B(n18), .C(n19), .D(n20), .Y(n2) );
  NAND4X1 U17 ( .A(n21), .B(n22), .C(n23), .D(n24), .Y(n20) );
  XNOR2X1 U18 ( .A(B[20]), .B(A[20]), .Y(n24) );
  XNOR2X1 U19 ( .A(B[21]), .B(A[21]), .Y(n23) );
  XNOR2X1 U20 ( .A(B[22]), .B(A[22]), .Y(n22) );
  XNOR2X1 U21 ( .A(B[23]), .B(A[23]), .Y(n21) );
  NAND4X1 U22 ( .A(n25), .B(n26), .C(n27), .D(n28), .Y(n19) );
  XNOR2X1 U23 ( .A(B[16]), .B(A[16]), .Y(n28) );
  XNOR2X1 U24 ( .A(B[17]), .B(A[17]), .Y(n27) );
  XNOR2X1 U25 ( .A(B[18]), .B(A[18]), .Y(n26) );
  XNOR2X1 U26 ( .A(B[19]), .B(A[19]), .Y(n25) );
  NAND4X1 U27 ( .A(n29), .B(n30), .C(n31), .D(n32), .Y(n18) );
  XNOR2X1 U28 ( .A(B[28]), .B(A[28]), .Y(n32) );
  XNOR2X1 U29 ( .A(B[29]), .B(A[29]), .Y(n31) );
  XNOR2X1 U30 ( .A(B[30]), .B(A[30]), .Y(n30) );
  XNOR2X1 U31 ( .A(B[31]), .B(A[31]), .Y(n29) );
  NAND4X1 U32 ( .A(n33), .B(n34), .C(n35), .D(n36), .Y(n17) );
  XNOR2X1 U33 ( .A(B[24]), .B(A[24]), .Y(n36) );
  XNOR2X1 U34 ( .A(B[25]), .B(A[25]), .Y(n35) );
  XNOR2X1 U35 ( .A(B[26]), .B(A[26]), .Y(n34) );
  XNOR2X1 U36 ( .A(B[27]), .B(A[27]), .Y(n33) );
  NOR2X1 U37 ( .A(n37), .B(n38), .Y(n1) );
  NAND4X1 U38 ( .A(n39), .B(n40), .C(n41), .D(n42), .Y(n38) );
  XNOR2X1 U39 ( .A(B[12]), .B(A[12]), .Y(n42) );
  XNOR2X1 U40 ( .A(B[13]), .B(A[13]), .Y(n41) );
  XNOR2X1 U41 ( .A(B[14]), .B(A[14]), .Y(n40) );
  XNOR2X1 U42 ( .A(B[15]), .B(A[15]), .Y(n39) );
  NAND4X1 U43 ( .A(n43), .B(n44), .C(n45), .D(n46), .Y(n37) );
  XNOR2X1 U44 ( .A(B[8]), .B(A[8]), .Y(n46) );
  XNOR2X1 U45 ( .A(B[9]), .B(A[9]), .Y(n45) );
  XNOR2X1 U46 ( .A(B[10]), .B(A[10]), .Y(n44) );
  XNOR2X1 U47 ( .A(B[11]), .B(A[11]), .Y(n43) );
endmodule


module CPU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[31] , \carry[30] , \carry[29] , \carry[28] ,
         \carry[27] , \carry[26] , \carry[25] , \carry[24] , \carry[23] ,
         \carry[22] , \carry[21] , \carry[20] , \carry[19] , \carry[18] ,
         \carry[17] , \carry[16] , \carry[15] , \carry[14] , \carry[13] ,
         \carry[12] , \carry[11] , \carry[10] , \carry[9] , \carry[8] ,
         \carry[7] , \carry[6] , \carry[5] , \carry[4] , \carry[3] ;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2X1 U1 ( .A(A[31]), .B(\carry[31] ), .Y(SUM[31]) );
  AND2X1 U2 ( .A(\carry[30] ), .B(A[30]), .Y(\carry[31] ) );
  XOR2X1 U3 ( .A(A[30]), .B(\carry[30] ), .Y(SUM[30]) );
  AND2X1 U4 ( .A(\carry[29] ), .B(A[29]), .Y(\carry[30] ) );
  XOR2X1 U5 ( .A(A[29]), .B(\carry[29] ), .Y(SUM[29]) );
  AND2X1 U6 ( .A(\carry[28] ), .B(A[28]), .Y(\carry[29] ) );
  XOR2X1 U7 ( .A(A[28]), .B(\carry[28] ), .Y(SUM[28]) );
  AND2X1 U8 ( .A(\carry[27] ), .B(A[27]), .Y(\carry[28] ) );
  XOR2X1 U9 ( .A(A[27]), .B(\carry[27] ), .Y(SUM[27]) );
  AND2X1 U10 ( .A(\carry[26] ), .B(A[26]), .Y(\carry[27] ) );
  XOR2X1 U11 ( .A(A[26]), .B(\carry[26] ), .Y(SUM[26]) );
  AND2X1 U12 ( .A(\carry[25] ), .B(A[25]), .Y(\carry[26] ) );
  XOR2X1 U13 ( .A(A[25]), .B(\carry[25] ), .Y(SUM[25]) );
  AND2X1 U14 ( .A(\carry[24] ), .B(A[24]), .Y(\carry[25] ) );
  XOR2X1 U15 ( .A(A[24]), .B(\carry[24] ), .Y(SUM[24]) );
  AND2X1 U16 ( .A(\carry[23] ), .B(A[23]), .Y(\carry[24] ) );
  XOR2X1 U17 ( .A(A[23]), .B(\carry[23] ), .Y(SUM[23]) );
  AND2X1 U18 ( .A(\carry[22] ), .B(A[22]), .Y(\carry[23] ) );
  XOR2X1 U19 ( .A(A[22]), .B(\carry[22] ), .Y(SUM[22]) );
  AND2X1 U20 ( .A(\carry[21] ), .B(A[21]), .Y(\carry[22] ) );
  XOR2X1 U21 ( .A(A[21]), .B(\carry[21] ), .Y(SUM[21]) );
  AND2X1 U22 ( .A(\carry[20] ), .B(A[20]), .Y(\carry[21] ) );
  XOR2X1 U23 ( .A(A[20]), .B(\carry[20] ), .Y(SUM[20]) );
  AND2X1 U24 ( .A(\carry[19] ), .B(A[19]), .Y(\carry[20] ) );
  XOR2X1 U25 ( .A(A[19]), .B(\carry[19] ), .Y(SUM[19]) );
  AND2X1 U26 ( .A(\carry[18] ), .B(A[18]), .Y(\carry[19] ) );
  XOR2X1 U27 ( .A(A[18]), .B(\carry[18] ), .Y(SUM[18]) );
  AND2X1 U28 ( .A(\carry[17] ), .B(A[17]), .Y(\carry[18] ) );
  XOR2X1 U29 ( .A(A[17]), .B(\carry[17] ), .Y(SUM[17]) );
  AND2X1 U30 ( .A(\carry[16] ), .B(A[16]), .Y(\carry[17] ) );
  XOR2X1 U31 ( .A(A[16]), .B(\carry[16] ), .Y(SUM[16]) );
  AND2X1 U32 ( .A(\carry[15] ), .B(A[15]), .Y(\carry[16] ) );
  XOR2X1 U33 ( .A(A[15]), .B(\carry[15] ), .Y(SUM[15]) );
  AND2X1 U34 ( .A(\carry[14] ), .B(A[14]), .Y(\carry[15] ) );
  XOR2X1 U35 ( .A(A[14]), .B(\carry[14] ), .Y(SUM[14]) );
  AND2X1 U36 ( .A(\carry[13] ), .B(A[13]), .Y(\carry[14] ) );
  XOR2X1 U37 ( .A(A[13]), .B(\carry[13] ), .Y(SUM[13]) );
  AND2X1 U38 ( .A(\carry[12] ), .B(A[12]), .Y(\carry[13] ) );
  XOR2X1 U39 ( .A(A[12]), .B(\carry[12] ), .Y(SUM[12]) );
  AND2X1 U40 ( .A(\carry[11] ), .B(A[11]), .Y(\carry[12] ) );
  XOR2X1 U41 ( .A(A[11]), .B(\carry[11] ), .Y(SUM[11]) );
  AND2X1 U42 ( .A(\carry[10] ), .B(A[10]), .Y(\carry[11] ) );
  XOR2X1 U43 ( .A(A[10]), .B(\carry[10] ), .Y(SUM[10]) );
  AND2X1 U44 ( .A(\carry[9] ), .B(A[9]), .Y(\carry[10] ) );
  XOR2X1 U45 ( .A(A[9]), .B(\carry[9] ), .Y(SUM[9]) );
  AND2X1 U46 ( .A(\carry[8] ), .B(A[8]), .Y(\carry[9] ) );
  XOR2X1 U47 ( .A(A[8]), .B(\carry[8] ), .Y(SUM[8]) );
  AND2X1 U48 ( .A(\carry[7] ), .B(A[7]), .Y(\carry[8] ) );
  XOR2X1 U49 ( .A(A[7]), .B(\carry[7] ), .Y(SUM[7]) );
  AND2X1 U50 ( .A(\carry[6] ), .B(A[6]), .Y(\carry[7] ) );
  XOR2X1 U51 ( .A(A[6]), .B(\carry[6] ), .Y(SUM[6]) );
  AND2X1 U52 ( .A(\carry[5] ), .B(A[5]), .Y(\carry[6] ) );
  XOR2X1 U53 ( .A(A[5]), .B(\carry[5] ), .Y(SUM[5]) );
  AND2X1 U54 ( .A(\carry[4] ), .B(A[4]), .Y(\carry[5] ) );
  XOR2X1 U55 ( .A(A[4]), .B(\carry[4] ), .Y(SUM[4]) );
  AND2X1 U56 ( .A(\carry[3] ), .B(A[3]), .Y(\carry[4] ) );
  XOR2X1 U57 ( .A(A[3]), .B(\carry[3] ), .Y(SUM[3]) );
  INVX1 U58 ( .A(\carry[3] ), .Y(SUM[2]) );
endmodule


module CPU_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] ;

  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        SUM[8]) );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        SUM[7]) );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        SUM[6]) );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        SUM[5]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(\carry[31] ), .Y(SUM[31]) );
  AND2X1 U1 ( .A(A[0]), .B(B[0]), .Y(\carry[1] ) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module detection ( stall, ena_data_out, addr_dst_out, addr1, addr2 );
  input [4:0] addr_dst_out;
  input [4:0] addr1;
  input [4:0] addr2;
  input ena_data_out;
  output stall;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  NOR2BX1 U1 ( .AN(ena_data_out), .B(n1), .Y(stall) );
  AOI33X1 U2 ( .A0(n2), .A1(n3), .A2(n4), .B0(n5), .B1(n6), .B2(n7), .Y(n1) );
  NOR3X1 U3 ( .A(n8), .B(n9), .C(n10), .Y(n7) );
  XOR2X1 U4 ( .A(addr_dst_out[3]), .B(addr1[3]), .Y(n10) );
  XOR2X1 U5 ( .A(addr_dst_out[1]), .B(addr1[1]), .Y(n9) );
  XOR2X1 U6 ( .A(addr_dst_out[0]), .B(addr1[0]), .Y(n8) );
  XNOR2X1 U7 ( .A(addr_dst_out[2]), .B(addr1[2]), .Y(n6) );
  XNOR2X1 U8 ( .A(addr_dst_out[4]), .B(addr1[4]), .Y(n5) );
  NOR3X1 U9 ( .A(n11), .B(n12), .C(n13), .Y(n4) );
  XOR2X1 U10 ( .A(addr_dst_out[3]), .B(addr2[3]), .Y(n13) );
  XOR2X1 U11 ( .A(addr_dst_out[1]), .B(addr2[1]), .Y(n12) );
  XOR2X1 U12 ( .A(addr_dst_out[0]), .B(addr2[0]), .Y(n11) );
  XNOR2X1 U13 ( .A(addr_dst_out[2]), .B(addr2[2]), .Y(n3) );
  XNOR2X1 U14 ( .A(addr_dst_out[4]), .B(addr2[4]), .Y(n2) );
endmodule


module Forward ( forwardA, forwardB, addr2_out, addr1_out, addr_dst_reg_out, 
        addr_dst_reg2_out, reg_rw_out_exe, reg_rw_out_mem, data_rw_reg_out, 
        sel_data_in, addr_dst, addr1, branch_ena, sel_data1, sel_data3, 
        addr_dst_out, addr2, sel_data2_in, sel_data1_in );
  output [1:0] forwardA;
  output [1:0] forwardB;
  input [4:0] addr2_out;
  input [4:0] addr1_out;
  input [4:0] addr_dst_reg_out;
  input [4:0] addr_dst_reg2_out;
  input [4:0] addr_dst;
  input [4:0] addr1;
  output [1:0] sel_data1;
  output [1:0] sel_data3;
  input [4:0] addr_dst_out;
  input [4:0] addr2;
  input reg_rw_out_exe, reg_rw_out_mem, data_rw_reg_out, branch_ena;
  output sel_data_in, sel_data2_in, sel_data1_in;
  wire   N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88;
  assign forwardA[1] = N33;

  NOR4X1 U1 ( .A(n1), .B(n2), .C(n3), .D(n4), .Y(sel_data_in) );
  XOR2X1 U2 ( .A(addr_dst_reg_out[1]), .B(addr_dst_reg2_out[1]), .Y(n4) );
  XOR2X1 U3 ( .A(addr_dst_reg_out[4]), .B(addr_dst_reg2_out[4]), .Y(n3) );
  XOR2X1 U4 ( .A(addr_dst_reg_out[2]), .B(addr_dst_reg2_out[2]), .Y(n2) );
  NAND3X1 U5 ( .A(n5), .B(data_rw_reg_out), .C(n6), .Y(n1) );
  XNOR2X1 U6 ( .A(addr_dst_reg_out[3]), .B(addr_dst_reg2_out[3]), .Y(n6) );
  XNOR2X1 U7 ( .A(addr_dst_reg_out[0]), .B(addr_dst_reg2_out[0]), .Y(n5) );
  NOR2X1 U8 ( .A(n7), .B(n8), .Y(sel_data3[1]) );
  AOI21X1 U9 ( .A0(branch_ena), .A1(n9), .B0(n10), .Y(n8) );
  INVX1 U10 ( .A(n11), .Y(n10) );
  NOR2X1 U11 ( .A(n12), .B(n13), .Y(sel_data3[0]) );
  AOI21X1 U12 ( .A0(n9), .A1(n11), .B0(n7), .Y(n12) );
  AND4X1 U13 ( .A(n14), .B(n15), .C(n16), .D(n17), .Y(n7) );
  NOR2X1 U14 ( .A(n18), .B(n19), .Y(n17) );
  XOR2X1 U15 ( .A(addr_dst_out[4]), .B(addr_dst[4]), .Y(n19) );
  XOR2X1 U16 ( .A(addr_dst_out[2]), .B(addr_dst[2]), .Y(n18) );
  XNOR2X1 U17 ( .A(addr_dst[0]), .B(addr_dst_out[0]), .Y(n16) );
  XNOR2X1 U18 ( .A(addr_dst[1]), .B(addr_dst_out[1]), .Y(n15) );
  XNOR2X1 U19 ( .A(addr_dst[3]), .B(addr_dst_out[3]), .Y(n14) );
  NAND4X1 U20 ( .A(n20), .B(n21), .C(n22), .D(n23), .Y(n11) );
  NOR3X1 U21 ( .A(n24), .B(n13), .C(n25), .Y(n23) );
  XOR2X1 U22 ( .A(addr_dst_reg_out[1]), .B(addr_dst[1]), .Y(n25) );
  XOR2X1 U23 ( .A(addr_dst_reg_out[0]), .B(addr_dst[0]), .Y(n24) );
  XNOR2X1 U24 ( .A(addr_dst[3]), .B(addr_dst_reg_out[3]), .Y(n22) );
  XNOR2X1 U25 ( .A(addr_dst[4]), .B(addr_dst_reg_out[4]), .Y(n21) );
  XNOR2X1 U26 ( .A(addr_dst[2]), .B(addr_dst_reg_out[2]), .Y(n20) );
  AND4X1 U27 ( .A(n26), .B(n27), .C(n28), .D(n29), .Y(n9) );
  NOR2X1 U28 ( .A(n30), .B(n31), .Y(n29) );
  XOR2X1 U29 ( .A(addr_dst_reg2_out[4]), .B(addr_dst[4]), .Y(n31) );
  XOR2X1 U30 ( .A(addr_dst_reg2_out[2]), .B(addr_dst[2]), .Y(n30) );
  XNOR2X1 U31 ( .A(addr_dst[0]), .B(addr_dst_reg2_out[0]), .Y(n28) );
  XNOR2X1 U32 ( .A(addr_dst[1]), .B(addr_dst_reg2_out[1]), .Y(n27) );
  XNOR2X1 U33 ( .A(addr_dst[3]), .B(addr_dst_reg2_out[3]), .Y(n26) );
  NOR4X1 U34 ( .A(n32), .B(n33), .C(n34), .D(n35), .Y(sel_data2_in) );
  XOR2X1 U35 ( .A(addr_dst_reg2_out[1]), .B(addr2[1]), .Y(n35) );
  XOR2X1 U36 ( .A(addr_dst_reg2_out[4]), .B(addr2[4]), .Y(n34) );
  XOR2X1 U37 ( .A(addr_dst_reg2_out[2]), .B(addr2[2]), .Y(n33) );
  NAND3X1 U38 ( .A(n36), .B(reg_rw_out_mem), .C(n37), .Y(n32) );
  XNOR2X1 U39 ( .A(addr_dst_reg2_out[3]), .B(addr2[3]), .Y(n37) );
  XNOR2X1 U40 ( .A(addr_dst_reg2_out[0]), .B(addr2[0]), .Y(n36) );
  NOR2BX1 U41 ( .AN(reg_rw_out_mem), .B(n38), .Y(sel_data1_in) );
  NOR2BX1 U42 ( .AN(n39), .B(n40), .Y(sel_data1[1]) );
  OAI21XL U43 ( .A0(n38), .A1(n13), .B0(n41), .Y(n39) );
  NOR2X1 U44 ( .A(n42), .B(n13), .Y(sel_data1[0]) );
  AOI21X1 U45 ( .A0(n43), .A1(n41), .B0(n40), .Y(n42) );
  AND4X1 U46 ( .A(n44), .B(n45), .C(n46), .D(n47), .Y(n40) );
  NOR2X1 U47 ( .A(n48), .B(n49), .Y(n47) );
  XOR2X1 U48 ( .A(addr_dst_out[4]), .B(addr1[4]), .Y(n49) );
  XOR2X1 U49 ( .A(addr_dst_out[2]), .B(addr1[2]), .Y(n48) );
  XNOR2X1 U50 ( .A(addr1[0]), .B(addr_dst_out[0]), .Y(n46) );
  XNOR2X1 U51 ( .A(addr1[1]), .B(addr_dst_out[1]), .Y(n45) );
  XNOR2X1 U52 ( .A(addr1[3]), .B(addr_dst_out[3]), .Y(n44) );
  NAND4X1 U53 ( .A(n50), .B(n51), .C(n52), .D(n53), .Y(n41) );
  NOR3X1 U54 ( .A(n54), .B(n13), .C(n55), .Y(n53) );
  XOR2X1 U55 ( .A(addr_dst_reg_out[1]), .B(addr1[1]), .Y(n55) );
  INVX1 U56 ( .A(branch_ena), .Y(n13) );
  XOR2X1 U57 ( .A(addr_dst_reg_out[0]), .B(addr1[0]), .Y(n54) );
  XNOR2X1 U58 ( .A(addr1[3]), .B(addr_dst_reg_out[3]), .Y(n52) );
  XNOR2X1 U59 ( .A(addr1[4]), .B(addr_dst_reg_out[4]), .Y(n51) );
  XNOR2X1 U60 ( .A(addr1[2]), .B(addr_dst_reg_out[2]), .Y(n50) );
  INVX1 U61 ( .A(n38), .Y(n43) );
  NAND4X1 U62 ( .A(n56), .B(n57), .C(n58), .D(n59), .Y(n38) );
  NOR2X1 U63 ( .A(n60), .B(n61), .Y(n59) );
  XOR2X1 U64 ( .A(addr_dst_reg2_out[4]), .B(addr1[4]), .Y(n61) );
  XOR2X1 U65 ( .A(addr_dst_reg2_out[2]), .B(addr1[2]), .Y(n60) );
  XNOR2X1 U66 ( .A(addr1[0]), .B(addr_dst_reg2_out[0]), .Y(n58) );
  XNOR2X1 U67 ( .A(addr1[1]), .B(addr_dst_reg2_out[1]), .Y(n57) );
  XNOR2X1 U68 ( .A(addr1[3]), .B(addr_dst_reg2_out[3]), .Y(n56) );
  NOR4X1 U69 ( .A(n62), .B(n63), .C(n64), .D(n65), .Y(forwardB[1]) );
  XOR2X1 U70 ( .A(addr_dst_reg2_out[1]), .B(addr2_out[1]), .Y(n65) );
  XOR2X1 U71 ( .A(addr_dst_reg2_out[4]), .B(addr2_out[4]), .Y(n64) );
  XOR2X1 U72 ( .A(addr_dst_reg2_out[2]), .B(addr2_out[2]), .Y(n63) );
  NAND4X1 U73 ( .A(n66), .B(n67), .C(reg_rw_out_mem), .D(n68), .Y(n62) );
  XNOR2X1 U74 ( .A(addr2_out[3]), .B(addr_dst_reg2_out[3]), .Y(n67) );
  XNOR2X1 U75 ( .A(addr2_out[0]), .B(addr_dst_reg2_out[0]), .Y(n66) );
  INVX1 U76 ( .A(n68), .Y(forwardB[0]) );
  NAND4X1 U77 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(n68) );
  NOR3X1 U78 ( .A(n73), .B(n74), .C(n75), .Y(n72) );
  XOR2X1 U79 ( .A(addr_dst_reg_out[1]), .B(addr2_out[1]), .Y(n75) );
  XOR2X1 U80 ( .A(addr_dst_reg_out[0]), .B(addr2_out[0]), .Y(n73) );
  XNOR2X1 U81 ( .A(addr2_out[3]), .B(addr_dst_reg_out[3]), .Y(n71) );
  XNOR2X1 U82 ( .A(addr2_out[4]), .B(addr_dst_reg_out[4]), .Y(n70) );
  XNOR2X1 U83 ( .A(addr2_out[2]), .B(addr_dst_reg_out[2]), .Y(n69) );
  INVX1 U84 ( .A(n76), .Y(forwardA[0]) );
  NOR4X1 U85 ( .A(n77), .B(n78), .C(n79), .D(n80), .Y(N33) );
  XOR2X1 U86 ( .A(addr_dst_reg2_out[1]), .B(addr1_out[1]), .Y(n80) );
  XOR2X1 U87 ( .A(addr_dst_reg2_out[4]), .B(addr1_out[4]), .Y(n79) );
  XOR2X1 U88 ( .A(addr_dst_reg2_out[2]), .B(addr1_out[2]), .Y(n78) );
  NAND4X1 U89 ( .A(n81), .B(n82), .C(reg_rw_out_mem), .D(n76), .Y(n77) );
  NAND4X1 U90 ( .A(n83), .B(n84), .C(n85), .D(n86), .Y(n76) );
  NOR3X1 U91 ( .A(n87), .B(n74), .C(n88), .Y(n86) );
  XOR2X1 U92 ( .A(addr_dst_reg_out[1]), .B(addr1_out[1]), .Y(n88) );
  INVX1 U93 ( .A(reg_rw_out_exe), .Y(n74) );
  XOR2X1 U94 ( .A(addr_dst_reg_out[0]), .B(addr1_out[0]), .Y(n87) );
  XNOR2X1 U95 ( .A(addr1_out[3]), .B(addr_dst_reg_out[3]), .Y(n85) );
  XNOR2X1 U96 ( .A(addr1_out[4]), .B(addr_dst_reg_out[4]), .Y(n84) );
  XNOR2X1 U97 ( .A(addr1_out[2]), .B(addr_dst_reg_out[2]), .Y(n83) );
  XNOR2X1 U98 ( .A(addr1_out[3]), .B(addr_dst_reg2_out[3]), .Y(n82) );
  XNOR2X1 U99 ( .A(addr1_out[0]), .B(addr_dst_reg2_out[0]), .Y(n81) );
endmodule


module MEMWB ( sel_wb_out, reg_rw_out, addr_dst_out, alu_result_out, 
        data_out_out, alu_result_in, sel_wb_in, reg_rw_in, addr_dst_in, 
        data_out_in, clk, rst );
  output [4:0] addr_dst_out;
  output [31:0] alu_result_out;
  output [31:0] data_out_out;
  input [31:0] alu_result_in;
  input [4:0] addr_dst_in;
  input [31:0] data_out_in;
  input sel_wb_in, reg_rw_in, clk, rst;
  output sel_wb_out, reg_rw_out;


  DFFRHQX1 \data_out_out_reg[31]  ( .D(data_out_in[31]), .CK(clk), .RN(rst), 
        .Q(data_out_out[31]) );
  DFFRHQX1 \data_out_out_reg[30]  ( .D(data_out_in[30]), .CK(clk), .RN(rst), 
        .Q(data_out_out[30]) );
  DFFRHQX1 \data_out_out_reg[29]  ( .D(data_out_in[29]), .CK(clk), .RN(rst), 
        .Q(data_out_out[29]) );
  DFFRHQX1 \data_out_out_reg[28]  ( .D(data_out_in[28]), .CK(clk), .RN(rst), 
        .Q(data_out_out[28]) );
  DFFRHQX1 \data_out_out_reg[27]  ( .D(data_out_in[27]), .CK(clk), .RN(rst), 
        .Q(data_out_out[27]) );
  DFFRHQX1 \data_out_out_reg[26]  ( .D(data_out_in[26]), .CK(clk), .RN(rst), 
        .Q(data_out_out[26]) );
  DFFRHQX1 \data_out_out_reg[25]  ( .D(data_out_in[25]), .CK(clk), .RN(rst), 
        .Q(data_out_out[25]) );
  DFFRHQX1 \data_out_out_reg[24]  ( .D(data_out_in[24]), .CK(clk), .RN(rst), 
        .Q(data_out_out[24]) );
  DFFRHQX1 \data_out_out_reg[23]  ( .D(data_out_in[23]), .CK(clk), .RN(rst), 
        .Q(data_out_out[23]) );
  DFFRHQX1 \data_out_out_reg[22]  ( .D(data_out_in[22]), .CK(clk), .RN(rst), 
        .Q(data_out_out[22]) );
  DFFRHQX1 \data_out_out_reg[21]  ( .D(data_out_in[21]), .CK(clk), .RN(rst), 
        .Q(data_out_out[21]) );
  DFFRHQX1 \data_out_out_reg[20]  ( .D(data_out_in[20]), .CK(clk), .RN(rst), 
        .Q(data_out_out[20]) );
  DFFRHQX1 \data_out_out_reg[19]  ( .D(data_out_in[19]), .CK(clk), .RN(rst), 
        .Q(data_out_out[19]) );
  DFFRHQX1 \data_out_out_reg[18]  ( .D(data_out_in[18]), .CK(clk), .RN(rst), 
        .Q(data_out_out[18]) );
  DFFRHQX1 \data_out_out_reg[17]  ( .D(data_out_in[17]), .CK(clk), .RN(rst), 
        .Q(data_out_out[17]) );
  DFFRHQX1 \data_out_out_reg[16]  ( .D(data_out_in[16]), .CK(clk), .RN(rst), 
        .Q(data_out_out[16]) );
  DFFRHQX1 \data_out_out_reg[15]  ( .D(data_out_in[15]), .CK(clk), .RN(rst), 
        .Q(data_out_out[15]) );
  DFFRHQX1 \alu_result_out_reg[31]  ( .D(alu_result_in[31]), .CK(clk), .RN(rst), .Q(alu_result_out[31]) );
  DFFRHQX1 \alu_result_out_reg[30]  ( .D(alu_result_in[30]), .CK(clk), .RN(rst), .Q(alu_result_out[30]) );
  DFFRHQX1 \alu_result_out_reg[29]  ( .D(alu_result_in[29]), .CK(clk), .RN(rst), .Q(alu_result_out[29]) );
  DFFRHQX1 \alu_result_out_reg[28]  ( .D(alu_result_in[28]), .CK(clk), .RN(rst), .Q(alu_result_out[28]) );
  DFFRHQX1 \alu_result_out_reg[27]  ( .D(alu_result_in[27]), .CK(clk), .RN(rst), .Q(alu_result_out[27]) );
  DFFRHQX1 \alu_result_out_reg[26]  ( .D(alu_result_in[26]), .CK(clk), .RN(rst), .Q(alu_result_out[26]) );
  DFFRHQX1 \alu_result_out_reg[25]  ( .D(alu_result_in[25]), .CK(clk), .RN(rst), .Q(alu_result_out[25]) );
  DFFRHQX1 \alu_result_out_reg[24]  ( .D(alu_result_in[24]), .CK(clk), .RN(rst), .Q(alu_result_out[24]) );
  DFFRHQX1 \alu_result_out_reg[23]  ( .D(alu_result_in[23]), .CK(clk), .RN(rst), .Q(alu_result_out[23]) );
  DFFRHQX1 \alu_result_out_reg[22]  ( .D(alu_result_in[22]), .CK(clk), .RN(rst), .Q(alu_result_out[22]) );
  DFFRHQX1 \alu_result_out_reg[21]  ( .D(alu_result_in[21]), .CK(clk), .RN(rst), .Q(alu_result_out[21]) );
  DFFRHQX1 \alu_result_out_reg[20]  ( .D(alu_result_in[20]), .CK(clk), .RN(rst), .Q(alu_result_out[20]) );
  DFFRHQX1 \alu_result_out_reg[19]  ( .D(alu_result_in[19]), .CK(clk), .RN(rst), .Q(alu_result_out[19]) );
  DFFRHQX1 \alu_result_out_reg[18]  ( .D(alu_result_in[18]), .CK(clk), .RN(rst), .Q(alu_result_out[18]) );
  DFFRHQX1 \alu_result_out_reg[17]  ( .D(alu_result_in[17]), .CK(clk), .RN(rst), .Q(alu_result_out[17]) );
  DFFRHQX1 \alu_result_out_reg[16]  ( .D(alu_result_in[16]), .CK(clk), .RN(rst), .Q(alu_result_out[16]) );
  DFFRHQX1 \alu_result_out_reg[15]  ( .D(alu_result_in[15]), .CK(clk), .RN(rst), .Q(alu_result_out[15]) );
  DFFRHQX1 \data_out_out_reg[14]  ( .D(data_out_in[14]), .CK(clk), .RN(rst), 
        .Q(data_out_out[14]) );
  DFFRHQX1 \data_out_out_reg[13]  ( .D(data_out_in[13]), .CK(clk), .RN(rst), 
        .Q(data_out_out[13]) );
  DFFRHQX1 \data_out_out_reg[12]  ( .D(data_out_in[12]), .CK(clk), .RN(rst), 
        .Q(data_out_out[12]) );
  DFFRHQX1 \data_out_out_reg[11]  ( .D(data_out_in[11]), .CK(clk), .RN(rst), 
        .Q(data_out_out[11]) );
  DFFRHQX1 \data_out_out_reg[10]  ( .D(data_out_in[10]), .CK(clk), .RN(rst), 
        .Q(data_out_out[10]) );
  DFFRHQX1 \data_out_out_reg[9]  ( .D(data_out_in[9]), .CK(clk), .RN(rst), .Q(
        data_out_out[9]) );
  DFFRHQX1 \data_out_out_reg[8]  ( .D(data_out_in[8]), .CK(clk), .RN(rst), .Q(
        data_out_out[8]) );
  DFFRHQX1 \data_out_out_reg[7]  ( .D(data_out_in[7]), .CK(clk), .RN(rst), .Q(
        data_out_out[7]) );
  DFFRHQX1 \data_out_out_reg[6]  ( .D(data_out_in[6]), .CK(clk), .RN(rst), .Q(
        data_out_out[6]) );
  DFFRHQX1 \data_out_out_reg[5]  ( .D(data_out_in[5]), .CK(clk), .RN(rst), .Q(
        data_out_out[5]) );
  DFFRHQX1 \data_out_out_reg[4]  ( .D(data_out_in[4]), .CK(clk), .RN(rst), .Q(
        data_out_out[4]) );
  DFFRHQX1 \data_out_out_reg[3]  ( .D(data_out_in[3]), .CK(clk), .RN(rst), .Q(
        data_out_out[3]) );
  DFFRHQX1 \alu_result_out_reg[14]  ( .D(alu_result_in[14]), .CK(clk), .RN(rst), .Q(alu_result_out[14]) );
  DFFRHQX1 \alu_result_out_reg[13]  ( .D(alu_result_in[13]), .CK(clk), .RN(rst), .Q(alu_result_out[13]) );
  DFFRHQX1 \alu_result_out_reg[12]  ( .D(alu_result_in[12]), .CK(clk), .RN(rst), .Q(alu_result_out[12]) );
  DFFRHQX1 \alu_result_out_reg[11]  ( .D(alu_result_in[11]), .CK(clk), .RN(rst), .Q(alu_result_out[11]) );
  DFFRHQX1 \alu_result_out_reg[10]  ( .D(alu_result_in[10]), .CK(clk), .RN(rst), .Q(alu_result_out[10]) );
  DFFRHQX1 \alu_result_out_reg[8]  ( .D(alu_result_in[8]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[8]) );
  DFFRHQX1 \alu_result_out_reg[7]  ( .D(alu_result_in[7]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[7]) );
  DFFRHQX1 \alu_result_out_reg[6]  ( .D(alu_result_in[6]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[6]) );
  DFFRHQX1 \alu_result_out_reg[5]  ( .D(alu_result_in[5]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[5]) );
  DFFRHQX1 \alu_result_out_reg[4]  ( .D(alu_result_in[4]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[4]) );
  DFFRHQX1 \alu_result_out_reg[3]  ( .D(alu_result_in[3]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[3]) );
  DFFRHQX1 \alu_result_out_reg[9]  ( .D(alu_result_in[9]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[9]) );
  DFFRHQX1 \data_out_out_reg[2]  ( .D(data_out_in[2]), .CK(clk), .RN(rst), .Q(
        data_out_out[2]) );
  DFFRHQX1 \data_out_out_reg[1]  ( .D(data_out_in[1]), .CK(clk), .RN(rst), .Q(
        data_out_out[1]) );
  DFFRHQX1 \data_out_out_reg[0]  ( .D(data_out_in[0]), .CK(clk), .RN(rst), .Q(
        data_out_out[0]) );
  DFFRHQX1 \alu_result_out_reg[2]  ( .D(alu_result_in[2]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[2]) );
  DFFRHQX1 \alu_result_out_reg[1]  ( .D(alu_result_in[1]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[1]) );
  DFFRHQX1 \alu_result_out_reg[0]  ( .D(alu_result_in[0]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[0]) );
  DFFRHQX1 reg_rw_out_reg ( .D(reg_rw_in), .CK(clk), .RN(rst), .Q(reg_rw_out)
         );
  DFFRHQX1 sel_wb_out_reg ( .D(sel_wb_in), .CK(clk), .RN(rst), .Q(sel_wb_out)
         );
  DFFRHQX1 \addr_dst_out_reg[4]  ( .D(addr_dst_in[4]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[4]) );
  DFFRHQX1 \addr_dst_out_reg[1]  ( .D(addr_dst_in[1]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[1]) );
  DFFRHQX1 \addr_dst_out_reg[2]  ( .D(addr_dst_in[2]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[2]) );
  DFFRHQX1 \addr_dst_out_reg[3]  ( .D(addr_dst_in[3]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[3]) );
  DFFRHQX1 \addr_dst_out_reg[0]  ( .D(addr_dst_in[0]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[0]) );
endmodule


module EXMEM ( ena_data_out, data_rw_out, sel_wb_out, reg_rw_out, 
        alu_result_out, read_data3_out, addr_dst_out, ena_data_in, data_rw_in, 
        sel_wb_in, reg_rw_in, alu_result_in, read_data3_in, addr_dst_in, clk, 
        rst );
  output [31:0] alu_result_out;
  output [31:0] read_data3_out;
  output [4:0] addr_dst_out;
  input [31:0] alu_result_in;
  input [31:0] read_data3_in;
  input [4:0] addr_dst_in;
  input ena_data_in, data_rw_in, sel_wb_in, reg_rw_in, clk, rst;
  output ena_data_out, data_rw_out, sel_wb_out, reg_rw_out;


  DFFRHQX1 data_rw_out_reg ( .D(data_rw_in), .CK(clk), .RN(rst), .Q(
        data_rw_out) );
  DFFRHQX1 \read_data3_out_reg[31]  ( .D(read_data3_in[31]), .CK(clk), .RN(rst), .Q(read_data3_out[31]) );
  DFFRHQX1 \read_data3_out_reg[30]  ( .D(read_data3_in[30]), .CK(clk), .RN(rst), .Q(read_data3_out[30]) );
  DFFRHQX1 \read_data3_out_reg[29]  ( .D(read_data3_in[29]), .CK(clk), .RN(rst), .Q(read_data3_out[29]) );
  DFFRHQX1 \read_data3_out_reg[28]  ( .D(read_data3_in[28]), .CK(clk), .RN(rst), .Q(read_data3_out[28]) );
  DFFRHQX1 \read_data3_out_reg[27]  ( .D(read_data3_in[27]), .CK(clk), .RN(rst), .Q(read_data3_out[27]) );
  DFFRHQX1 \read_data3_out_reg[26]  ( .D(read_data3_in[26]), .CK(clk), .RN(rst), .Q(read_data3_out[26]) );
  DFFRHQX1 \read_data3_out_reg[25]  ( .D(read_data3_in[25]), .CK(clk), .RN(rst), .Q(read_data3_out[25]) );
  DFFRHQX1 \read_data3_out_reg[24]  ( .D(read_data3_in[24]), .CK(clk), .RN(rst), .Q(read_data3_out[24]) );
  DFFRHQX1 \read_data3_out_reg[23]  ( .D(read_data3_in[23]), .CK(clk), .RN(rst), .Q(read_data3_out[23]) );
  DFFRHQX1 \read_data3_out_reg[22]  ( .D(read_data3_in[22]), .CK(clk), .RN(rst), .Q(read_data3_out[22]) );
  DFFRHQX1 \read_data3_out_reg[21]  ( .D(read_data3_in[21]), .CK(clk), .RN(rst), .Q(read_data3_out[21]) );
  DFFRHQX1 \read_data3_out_reg[20]  ( .D(read_data3_in[20]), .CK(clk), .RN(rst), .Q(read_data3_out[20]) );
  DFFRHQX1 \read_data3_out_reg[19]  ( .D(read_data3_in[19]), .CK(clk), .RN(rst), .Q(read_data3_out[19]) );
  DFFRHQX1 \read_data3_out_reg[18]  ( .D(read_data3_in[18]), .CK(clk), .RN(rst), .Q(read_data3_out[18]) );
  DFFRHQX1 \read_data3_out_reg[17]  ( .D(read_data3_in[17]), .CK(clk), .RN(rst), .Q(read_data3_out[17]) );
  DFFRHQX1 \read_data3_out_reg[16]  ( .D(read_data3_in[16]), .CK(clk), .RN(rst), .Q(read_data3_out[16]) );
  DFFRHQX1 \read_data3_out_reg[15]  ( .D(read_data3_in[15]), .CK(clk), .RN(rst), .Q(read_data3_out[15]) );
  DFFRHQX1 \read_data3_out_reg[14]  ( .D(read_data3_in[14]), .CK(clk), .RN(rst), .Q(read_data3_out[14]) );
  DFFRHQX1 \read_data3_out_reg[13]  ( .D(read_data3_in[13]), .CK(clk), .RN(rst), .Q(read_data3_out[13]) );
  DFFRHQX1 \read_data3_out_reg[12]  ( .D(read_data3_in[12]), .CK(clk), .RN(rst), .Q(read_data3_out[12]) );
  DFFRHQX1 \read_data3_out_reg[11]  ( .D(read_data3_in[11]), .CK(clk), .RN(rst), .Q(read_data3_out[11]) );
  DFFRHQX1 \read_data3_out_reg[10]  ( .D(read_data3_in[10]), .CK(clk), .RN(rst), .Q(read_data3_out[10]) );
  DFFRHQX1 \read_data3_out_reg[9]  ( .D(read_data3_in[9]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[9]) );
  DFFRHQX1 \read_data3_out_reg[8]  ( .D(read_data3_in[8]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[8]) );
  DFFRHQX1 \read_data3_out_reg[7]  ( .D(read_data3_in[7]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[7]) );
  DFFRHQX1 \read_data3_out_reg[6]  ( .D(read_data3_in[6]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[6]) );
  DFFRHQX1 \read_data3_out_reg[5]  ( .D(read_data3_in[5]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[5]) );
  DFFRHQX1 \read_data3_out_reg[4]  ( .D(read_data3_in[4]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[4]) );
  DFFRHQX1 \read_data3_out_reg[3]  ( .D(read_data3_in[3]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[3]) );
  DFFRHQX1 \read_data3_out_reg[2]  ( .D(read_data3_in[2]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[2]) );
  DFFRHQX1 \read_data3_out_reg[1]  ( .D(read_data3_in[1]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[1]) );
  DFFRHQX1 \read_data3_out_reg[0]  ( .D(read_data3_in[0]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[0]) );
  DFFRHQX1 \alu_result_out_reg[31]  ( .D(alu_result_in[31]), .CK(clk), .RN(rst), .Q(alu_result_out[31]) );
  DFFRHQX1 \alu_result_out_reg[30]  ( .D(alu_result_in[30]), .CK(clk), .RN(rst), .Q(alu_result_out[30]) );
  DFFRHQX1 \alu_result_out_reg[29]  ( .D(alu_result_in[29]), .CK(clk), .RN(rst), .Q(alu_result_out[29]) );
  DFFRHQX1 \alu_result_out_reg[28]  ( .D(alu_result_in[28]), .CK(clk), .RN(rst), .Q(alu_result_out[28]) );
  DFFRHQX1 \alu_result_out_reg[27]  ( .D(alu_result_in[27]), .CK(clk), .RN(rst), .Q(alu_result_out[27]) );
  DFFRHQX1 \alu_result_out_reg[26]  ( .D(alu_result_in[26]), .CK(clk), .RN(rst), .Q(alu_result_out[26]) );
  DFFRHQX1 \alu_result_out_reg[25]  ( .D(alu_result_in[25]), .CK(clk), .RN(rst), .Q(alu_result_out[25]) );
  DFFRHQX1 \alu_result_out_reg[24]  ( .D(alu_result_in[24]), .CK(clk), .RN(rst), .Q(alu_result_out[24]) );
  DFFRHQX1 \alu_result_out_reg[23]  ( .D(alu_result_in[23]), .CK(clk), .RN(rst), .Q(alu_result_out[23]) );
  DFFRHQX1 \alu_result_out_reg[22]  ( .D(alu_result_in[22]), .CK(clk), .RN(rst), .Q(alu_result_out[22]) );
  DFFRHQX1 \alu_result_out_reg[21]  ( .D(alu_result_in[21]), .CK(clk), .RN(rst), .Q(alu_result_out[21]) );
  DFFRHQX1 \alu_result_out_reg[20]  ( .D(alu_result_in[20]), .CK(clk), .RN(rst), .Q(alu_result_out[20]) );
  DFFRHQX1 \alu_result_out_reg[19]  ( .D(alu_result_in[19]), .CK(clk), .RN(rst), .Q(alu_result_out[19]) );
  DFFRHQX1 \alu_result_out_reg[18]  ( .D(alu_result_in[18]), .CK(clk), .RN(rst), .Q(alu_result_out[18]) );
  DFFRHQX1 \alu_result_out_reg[17]  ( .D(alu_result_in[17]), .CK(clk), .RN(rst), .Q(alu_result_out[17]) );
  DFFRHQX1 \alu_result_out_reg[16]  ( .D(alu_result_in[16]), .CK(clk), .RN(rst), .Q(alu_result_out[16]) );
  DFFRHQX1 \alu_result_out_reg[15]  ( .D(alu_result_in[15]), .CK(clk), .RN(rst), .Q(alu_result_out[15]) );
  DFFRHQX1 \alu_result_out_reg[14]  ( .D(alu_result_in[14]), .CK(clk), .RN(rst), .Q(alu_result_out[14]) );
  DFFRHQX1 \alu_result_out_reg[13]  ( .D(alu_result_in[13]), .CK(clk), .RN(rst), .Q(alu_result_out[13]) );
  DFFRHQX1 \alu_result_out_reg[12]  ( .D(alu_result_in[12]), .CK(clk), .RN(rst), .Q(alu_result_out[12]) );
  DFFRHQX1 \alu_result_out_reg[11]  ( .D(alu_result_in[11]), .CK(clk), .RN(rst), .Q(alu_result_out[11]) );
  DFFRHQX1 \alu_result_out_reg[10]  ( .D(alu_result_in[10]), .CK(clk), .RN(rst), .Q(alu_result_out[10]) );
  DFFRHQX1 \alu_result_out_reg[9]  ( .D(alu_result_in[9]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[9]) );
  DFFRHQX1 \alu_result_out_reg[8]  ( .D(alu_result_in[8]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[8]) );
  DFFRHQX1 \alu_result_out_reg[7]  ( .D(alu_result_in[7]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[7]) );
  DFFRHQX1 \alu_result_out_reg[6]  ( .D(alu_result_in[6]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[6]) );
  DFFRHQX1 \alu_result_out_reg[5]  ( .D(alu_result_in[5]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[5]) );
  DFFRHQX1 \alu_result_out_reg[4]  ( .D(alu_result_in[4]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[4]) );
  DFFRHQX1 \alu_result_out_reg[3]  ( .D(alu_result_in[3]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[3]) );
  DFFRHQX1 reg_rw_out_reg ( .D(reg_rw_in), .CK(clk), .RN(rst), .Q(reg_rw_out)
         );
  DFFRHQX1 \alu_result_out_reg[2]  ( .D(alu_result_in[2]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[2]) );
  DFFRHQX1 \alu_result_out_reg[1]  ( .D(alu_result_in[1]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[1]) );
  DFFRHQX1 \alu_result_out_reg[0]  ( .D(alu_result_in[0]), .CK(clk), .RN(rst), 
        .Q(alu_result_out[0]) );
  DFFRHQX1 \addr_dst_out_reg[1]  ( .D(addr_dst_in[1]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[1]) );
  DFFRHQX1 \addr_dst_out_reg[0]  ( .D(addr_dst_in[0]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[0]) );
  DFFRHQX1 \addr_dst_out_reg[4]  ( .D(addr_dst_in[4]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[4]) );
  DFFRHQX1 \addr_dst_out_reg[2]  ( .D(addr_dst_in[2]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[2]) );
  DFFRHQX1 \addr_dst_out_reg[3]  ( .D(addr_dst_in[3]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[3]) );
  DFFRHQX1 ena_data_out_reg ( .D(ena_data_in), .CK(clk), .RN(rst), .Q(
        ena_data_out) );
  DFFRHQX1 sel_wb_out_reg ( .D(sel_wb_in), .CK(clk), .RN(rst), .Q(sel_wb_out)
         );
endmodule


module ALU ( ls_w_mode, funct, sv, source1, source2, over_flow, alu_result );
  input [3:0] funct;
  input [1:0] sv;
  input [31:0] source1;
  input [31:0] source2;
  output [31:0] alu_result;
  input ls_w_mode;
  output over_flow;
  wire   N14, N15, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, \offset[9] , \offset[8] , \offset[7] ,
         \offset[6] , \offset[5] , \offset[4] , \offset[3] , \offset[31] ,
         \offset[30] , \offset[2] , \offset[29] , \offset[28] , \offset[27] ,
         \offset[26] , \offset[25] , \offset[24] , \offset[23] , \offset[22] ,
         \offset[21] , \offset[20] , \offset[1] , \offset[19] , \offset[18] ,
         \offset[17] , \offset[16] , \offset[15] , \offset[14] , \offset[13] ,
         \offset[12] , \offset[11] , \offset[10] , \offset[0] , n64, n65, n66,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n84, n85, n87, n88,
         n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n101, n102, n103,
         n104, n105, n106, n108, n109, n110, n111, n112, n113, n115, n116,
         n117, n118, n119, n120, n122, n123, n124, n125, n126, n127, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n142, n143, n144, n145, n146, n147, n149, n150, n151, n152, n153,
         n154, n156, n157, n158, n159, n160, n161, n163, n164, n165, n166,
         n167, n168, n170, n171, n172, n173, n174, n175, n177, n178, n179,
         n180, n181, n182, n184, n185, n186, n187, n188, n189, n191, n192,
         n193, n194, n195, n196, n198, n199, n200, n201, n202, n203, n205,
         n206, n207, n208, n209, n210, n212, n213, n214, n215, n216, n217,
         n219, n220, n221, n222, n223, n224, n226, n227, n228, n229, n230,
         n231, n233, n234, n235, n236, n237, n238, n240, n241, n242, n243,
         n244, n245, n247, n248, n249, n250, n251, n252, n254, n255, n256,
         n257, n258, n259, n261, n262, n263, n264, n265, n266, n268, n269,
         n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n282,
         n283, n284, n285, n286, n287, n289, n290, n291, n292, n293, n294,
         n296, n297, n298, n299, n300, n301, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n67, n78, n79, n80, n81, n82, n83, n86, n93, n100,
         n107, n114, n121, n128, n141, n148, n155, n162, n169, n176, n183,
         n190, n197, n204, n211, n218, n225, n232, n239, n246, n253, n260,
         n267, n274, n281, n288, n295, n302, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508;
  wire   [31:0] rotate_tmp;

  ALU_DW01_add_0 add_79 ( .A({n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, 
        n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
        n34, n33, n32, n31, n30, n29, n28, n27}), .B({\offset[31] , 
        \offset[30] , \offset[29] , \offset[28] , \offset[27] , \offset[26] , 
        \offset[25] , \offset[24] , \offset[23] , \offset[22] , \offset[21] , 
        \offset[20] , \offset[19] , \offset[18] , \offset[17] , \offset[16] , 
        \offset[15] , \offset[14] , \offset[13] , \offset[12] , \offset[11] , 
        \offset[10] , \offset[9] , \offset[8] , \offset[7] , \offset[6] , 
        \offset[5] , \offset[4] , \offset[3] , \offset[2] , \offset[1] , 
        \offset[0] }), .CI(1'b0), .SUM({N284, N283, N282, N281, N280, N279, 
        N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, 
        N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, 
        N254, N253}) );
  ALU_DW01_ash_0 sll_74 ( .A({n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, 
        n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
        n34, n33, n32, n31, n30, n29, n28, n27}), .DATA_TC(1'b0), .SH({n26, 
        source2[30:6], n25, n24, n23, n21, n15, n14}), .SH_TC(1'b0), .B({N252, 
        N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, 
        N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, 
        N227, N226, N225, N224, N223, N222, N221}) );
  ALU_DW_rash_0 srl_64 ( .A({n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, 
        n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
        n34, n33, n32, n31, n30, n29, n28, n27}), .DATA_TC(1'b0), .SH({n26, 
        source2[30:6], n25, n24, n23, n21, n15, n14}), .SH_TC(1'b0), .B({N220, 
        N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, 
        N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, 
        N195, N194, N193, N192, N191, N190, N189}) );
  ALU_DW01_sub_0 sub_42 ( .A({n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, 
        n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
        n34, n33, n32, n31, n30, n29, n28, n27}), .B({n26, source2[30:6], n25, 
        n24, n23, n21, n15, n14}), .CI(1'b0), .DIFF({N285, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61}) );
  ALU_DW01_add_1 add_34 ( .A({n58, n57, n56, n55, n54, n53, n52, n51, n50, n49, 
        n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
        n34, n33, n32, n31, n30, n29, n28, n27}), .B({n26, source2[30:6], n25, 
        n24, n23, n21, n15, n14}), .CI(1'b0), .SUM({N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28}) );
  ALU_DW01_ash_1 sll_26 ( .A({n26, source2[30:6], n25, n24, n23, n21, n15, n14}), .DATA_TC(1'b0), .SH({N15, N14}), .SH_TC(1'b0), .B({\offset[31] , 
        \offset[30] , \offset[29] , \offset[28] , \offset[27] , \offset[26] , 
        \offset[25] , \offset[24] , \offset[23] , \offset[22] , \offset[21] , 
        \offset[20] , \offset[19] , \offset[18] , \offset[17] , \offset[16] , 
        \offset[15] , \offset[14] , \offset[13] , \offset[12] , \offset[11] , 
        \offset[10] , \offset[9] , \offset[8] , \offset[7] , \offset[6] , 
        \offset[5] , \offset[4] , \offset[3] , \offset[2] , \offset[1] , 
        \offset[0] }) );
  NOR2X1 U5 ( .A(n14), .B(n15), .Y(n1) );
  NAND3X1 U6 ( .A(n304), .B(n310), .C(funct[2]), .Y(n2) );
  NOR2X1 U7 ( .A(n21), .B(n23), .Y(n3) );
  NOR2X1 U8 ( .A(n107), .B(n302), .Y(n4) );
  NOR3X1 U9 ( .A(n307), .B(n311), .C(n309), .Y(n5) );
  OR3XL U10 ( .A(n306), .B(funct[1]), .C(n303), .Y(n6) );
  NOR2X1 U11 ( .A(n107), .B(n23), .Y(n7) );
  NOR2X1 U15 ( .A(n21), .B(n302), .Y(n8) );
  NOR3X1 U17 ( .A(n306), .B(funct[2]), .C(n310), .Y(n9) );
  NOR3X1 U18 ( .A(n310), .B(n306), .C(n303), .Y(n10) );
  NAND3X1 U19 ( .A(funct[1]), .B(n303), .C(n304), .Y(n11) );
  AND2X2 U20 ( .A(n86), .B(n15), .Y(n12) );
  NAND2X1 U21 ( .A(n358), .B(n24), .Y(n13) );
  INVX1 U22 ( .A(n336), .Y(n59) );
  INVX1 U23 ( .A(n331), .Y(n61) );
  INVX1 U24 ( .A(n12), .Y(n60) );
  INVX1 U25 ( .A(n305), .Y(n62) );
  AOI22X1 U26 ( .A0(N274), .A1(n5), .B0(N242), .B1(n84), .Y(n207) );
  AOI22X1 U27 ( .A0(N275), .A1(n5), .B0(N243), .B1(n84), .Y(n200) );
  AOI22X1 U28 ( .A0(N276), .A1(n5), .B0(N244), .B1(n84), .Y(n193) );
  AOI22X1 U29 ( .A0(N277), .A1(n5), .B0(N245), .B1(n84), .Y(n186) );
  AOI22X1 U30 ( .A0(N278), .A1(n5), .B0(N246), .B1(n84), .Y(n179) );
  AOI22X1 U31 ( .A0(N279), .A1(n5), .B0(N247), .B1(n84), .Y(n172) );
  AOI22X1 U32 ( .A0(N280), .A1(n5), .B0(N248), .B1(n84), .Y(n165) );
  AOI22X1 U33 ( .A0(N281), .A1(n5), .B0(N249), .B1(n84), .Y(n158) );
  AOI22X1 U34 ( .A0(N282), .A1(n5), .B0(N250), .B1(n84), .Y(n151) );
  AOI22X1 U35 ( .A0(N283), .A1(n5), .B0(N251), .B1(n84), .Y(n137) );
  AOI22X1 U36 ( .A0(N254), .A1(n5), .B0(N222), .B1(n84), .Y(n221) );
  AOI22X1 U37 ( .A0(N255), .A1(n5), .B0(N223), .B1(n84), .Y(n144) );
  AOI22X1 U38 ( .A0(N256), .A1(n5), .B0(N224), .B1(n84), .Y(n124) );
  AOI22X1 U39 ( .A0(N257), .A1(n5), .B0(N225), .B1(n84), .Y(n117) );
  AOI22X1 U40 ( .A0(N258), .A1(n5), .B0(N226), .B1(n84), .Y(n110) );
  AOI22X1 U41 ( .A0(N259), .A1(n5), .B0(N227), .B1(n84), .Y(n103) );
  AOI22X1 U42 ( .A0(N260), .A1(n5), .B0(N228), .B1(n84), .Y(n96) );
  AOI22X1 U43 ( .A0(N261), .A1(n5), .B0(N229), .B1(n84), .Y(n89) );
  AOI22X1 U44 ( .A0(N262), .A1(n5), .B0(N230), .B1(n84), .Y(n74) );
  AOI22X1 U45 ( .A0(N270), .A1(n5), .B0(N238), .B1(n84), .Y(n242) );
  AOI22X1 U46 ( .A0(N271), .A1(n5), .B0(N239), .B1(n84), .Y(n235) );
  AOI22X1 U47 ( .A0(N272), .A1(n5), .B0(N240), .B1(n84), .Y(n228) );
  AOI22X1 U48 ( .A0(N273), .A1(n5), .B0(N241), .B1(n84), .Y(n214) );
  AOI22X1 U49 ( .A0(N263), .A1(n5), .B0(N231), .B1(n84), .Y(n291) );
  AOI22X1 U50 ( .A0(N264), .A1(n5), .B0(N232), .B1(n84), .Y(n284) );
  AOI22X1 U51 ( .A0(N265), .A1(n5), .B0(N233), .B1(n84), .Y(n277) );
  AOI22X1 U52 ( .A0(N266), .A1(n5), .B0(N234), .B1(n84), .Y(n270) );
  AOI22X1 U53 ( .A0(N267), .A1(n5), .B0(N235), .B1(n84), .Y(n263) );
  AOI22X1 U54 ( .A0(N268), .A1(n5), .B0(N236), .B1(n84), .Y(n256) );
  AOI22X1 U55 ( .A0(N269), .A1(n5), .B0(N237), .B1(n84), .Y(n249) );
  NAND4X1 U56 ( .A(n156), .B(n157), .C(n158), .D(n159), .Y(alu_result[28]) );
  AOI22X1 U57 ( .A0(n55), .A1(n160), .B0(source2[28]), .B1(n161), .Y(n159) );
  AOI22X1 U58 ( .A0(rotate_tmp[28]), .A1(n85), .B0(N217), .B1(n10), .Y(n157)
         );
  AOI22X1 U59 ( .A0(N89), .A1(n9), .B0(N56), .B1(n69), .Y(n156) );
  NAND4X1 U60 ( .A(n170), .B(n171), .C(n172), .D(n173), .Y(alu_result[26]) );
  AOI22X1 U61 ( .A0(n53), .A1(n174), .B0(source2[26]), .B1(n175), .Y(n173) );
  AOI22X1 U62 ( .A0(rotate_tmp[26]), .A1(n85), .B0(N215), .B1(n10), .Y(n171)
         );
  AOI22X1 U63 ( .A0(N87), .A1(n9), .B0(N54), .B1(n69), .Y(n170) );
  NAND4X1 U64 ( .A(n163), .B(n164), .C(n165), .D(n166), .Y(alu_result[27]) );
  AOI22X1 U65 ( .A0(n54), .A1(n167), .B0(source2[27]), .B1(n168), .Y(n166) );
  AOI22X1 U66 ( .A0(rotate_tmp[27]), .A1(n85), .B0(N216), .B1(n10), .Y(n164)
         );
  AOI22X1 U67 ( .A0(N88), .A1(n9), .B0(N55), .B1(n69), .Y(n163) );
  NAND4X1 U68 ( .A(n198), .B(n199), .C(n200), .D(n201), .Y(alu_result[22]) );
  AOI22X1 U69 ( .A0(n49), .A1(n202), .B0(source2[22]), .B1(n203), .Y(n201) );
  AOI22X1 U70 ( .A0(rotate_tmp[22]), .A1(n85), .B0(N211), .B1(n10), .Y(n199)
         );
  AOI22X1 U71 ( .A0(N83), .A1(n9), .B0(N50), .B1(n69), .Y(n198) );
  NAND4X1 U72 ( .A(n177), .B(n178), .C(n179), .D(n180), .Y(alu_result[25]) );
  AOI22X1 U73 ( .A0(n52), .A1(n181), .B0(source2[25]), .B1(n182), .Y(n180) );
  AOI22X1 U74 ( .A0(rotate_tmp[25]), .A1(n85), .B0(N214), .B1(n10), .Y(n178)
         );
  AOI22X1 U75 ( .A0(N86), .A1(n9), .B0(N53), .B1(n69), .Y(n177) );
  NAND4X1 U76 ( .A(n149), .B(n150), .C(n151), .D(n152), .Y(alu_result[29]) );
  AOI22X1 U77 ( .A0(n56), .A1(n153), .B0(source2[29]), .B1(n154), .Y(n152) );
  AOI22X1 U78 ( .A0(rotate_tmp[29]), .A1(n85), .B0(N218), .B1(n10), .Y(n150)
         );
  AOI22X1 U79 ( .A0(N90), .A1(n9), .B0(N57), .B1(n69), .Y(n149) );
  NAND4X1 U80 ( .A(n184), .B(n185), .C(n186), .D(n187), .Y(alu_result[24]) );
  AOI22X1 U81 ( .A0(n51), .A1(n188), .B0(source2[24]), .B1(n189), .Y(n187) );
  AOI22X1 U82 ( .A0(rotate_tmp[24]), .A1(n85), .B0(N213), .B1(n10), .Y(n185)
         );
  AOI22X1 U83 ( .A0(N85), .A1(n9), .B0(N52), .B1(n69), .Y(n184) );
  NAND4X1 U84 ( .A(n135), .B(n136), .C(n137), .D(n138), .Y(alu_result[30]) );
  AOI22X1 U85 ( .A0(n57), .A1(n139), .B0(source2[30]), .B1(n140), .Y(n138) );
  AOI22X1 U86 ( .A0(rotate_tmp[30]), .A1(n85), .B0(N219), .B1(n10), .Y(n136)
         );
  AOI22X1 U87 ( .A0(N91), .A1(n9), .B0(N58), .B1(n69), .Y(n135) );
  NAND4X1 U88 ( .A(n191), .B(n192), .C(n193), .D(n194), .Y(alu_result[23]) );
  AOI22X1 U89 ( .A0(n50), .A1(n195), .B0(source2[23]), .B1(n196), .Y(n194) );
  AOI22X1 U90 ( .A0(rotate_tmp[23]), .A1(n85), .B0(N212), .B1(n10), .Y(n192)
         );
  AOI22X1 U91 ( .A0(N84), .A1(n9), .B0(N51), .B1(n69), .Y(n191) );
  NAND4X1 U92 ( .A(n205), .B(n206), .C(n207), .D(n208), .Y(alu_result[21]) );
  AOI22X1 U93 ( .A0(n48), .A1(n209), .B0(source2[21]), .B1(n210), .Y(n208) );
  AOI22X1 U94 ( .A0(rotate_tmp[21]), .A1(n85), .B0(N210), .B1(n10), .Y(n206)
         );
  AOI22X1 U95 ( .A0(N82), .A1(n9), .B0(N49), .B1(n69), .Y(n205) );
  NAND4X1 U96 ( .A(n129), .B(n130), .C(n131), .D(n132), .Y(alu_result[31]) );
  AOI22X1 U97 ( .A0(n58), .A1(n133), .B0(n26), .B1(n134), .Y(n132) );
  AOI22X1 U98 ( .A0(rotate_tmp[31]), .A1(n85), .B0(N220), .B1(n10), .Y(n130)
         );
  AOI22X1 U99 ( .A0(N285), .A1(n9), .B0(N59), .B1(n69), .Y(n129) );
  AOI22X1 U100 ( .A0(N284), .A1(n5), .B0(N252), .B1(n84), .Y(n131) );
  NAND4X1 U101 ( .A(n72), .B(n73), .C(n74), .D(n75), .Y(alu_result[9]) );
  AOI22X1 U102 ( .A0(n36), .A1(n76), .B0(source2[9]), .B1(n77), .Y(n75) );
  AOI22X1 U103 ( .A0(N70), .A1(n9), .B0(N37), .B1(n69), .Y(n72) );
  AOI22X1 U104 ( .A0(rotate_tmp[9]), .A1(n85), .B0(N198), .B1(n10), .Y(n73) );
  NAND4X1 U105 ( .A(n87), .B(n88), .C(n89), .D(n90), .Y(alu_result[8]) );
  AOI22X1 U106 ( .A0(n35), .A1(n91), .B0(source2[8]), .B1(n92), .Y(n90) );
  AOI22X1 U107 ( .A0(N69), .A1(n9), .B0(N36), .B1(n69), .Y(n87) );
  AOI22X1 U108 ( .A0(rotate_tmp[8]), .A1(n85), .B0(N197), .B1(n10), .Y(n88) );
  NAND4X1 U109 ( .A(n94), .B(n95), .C(n96), .D(n97), .Y(alu_result[7]) );
  AOI22X1 U110 ( .A0(n34), .A1(n98), .B0(source2[7]), .B1(n99), .Y(n97) );
  AOI22X1 U111 ( .A0(N68), .A1(n9), .B0(N35), .B1(n69), .Y(n94) );
  AOI22X1 U112 ( .A0(rotate_tmp[7]), .A1(n85), .B0(N196), .B1(n10), .Y(n95) );
  NAND4X1 U113 ( .A(n101), .B(n102), .C(n103), .D(n104), .Y(alu_result[6]) );
  AOI22X1 U114 ( .A0(n33), .A1(n105), .B0(source2[6]), .B1(n106), .Y(n104) );
  AOI22X1 U115 ( .A0(N67), .A1(n9), .B0(N34), .B1(n69), .Y(n101) );
  AOI22X1 U116 ( .A0(rotate_tmp[6]), .A1(n85), .B0(N195), .B1(n10), .Y(n102)
         );
  NAND4X1 U117 ( .A(n289), .B(n290), .C(n291), .D(n292), .Y(alu_result[10]) );
  AOI22X1 U118 ( .A0(n37), .A1(n293), .B0(source2[10]), .B1(n294), .Y(n292) );
  AOI22X1 U119 ( .A0(rotate_tmp[10]), .A1(n85), .B0(N199), .B1(n10), .Y(n290)
         );
  AOI22X1 U120 ( .A0(N71), .A1(n9), .B0(N38), .B1(n69), .Y(n289) );
  NAND4X1 U121 ( .A(n247), .B(n248), .C(n249), .D(n250), .Y(alu_result[16]) );
  AOI22X1 U122 ( .A0(n43), .A1(n251), .B0(source2[16]), .B1(n252), .Y(n250) );
  AOI22X1 U123 ( .A0(rotate_tmp[16]), .A1(n85), .B0(N205), .B1(n10), .Y(n248)
         );
  AOI22X1 U124 ( .A0(N77), .A1(n9), .B0(N44), .B1(n69), .Y(n247) );
  NAND4X1 U125 ( .A(n233), .B(n234), .C(n235), .D(n236), .Y(alu_result[18]) );
  AOI22X1 U126 ( .A0(n45), .A1(n237), .B0(source2[18]), .B1(n238), .Y(n236) );
  AOI22X1 U127 ( .A0(rotate_tmp[18]), .A1(n85), .B0(N207), .B1(n10), .Y(n234)
         );
  AOI22X1 U128 ( .A0(N79), .A1(n9), .B0(N46), .B1(n69), .Y(n233) );
  NAND4X1 U129 ( .A(n275), .B(n276), .C(n277), .D(n278), .Y(alu_result[12]) );
  AOI22X1 U130 ( .A0(n39), .A1(n279), .B0(source2[12]), .B1(n280), .Y(n278) );
  AOI22X1 U131 ( .A0(rotate_tmp[12]), .A1(n85), .B0(N201), .B1(n10), .Y(n276)
         );
  AOI22X1 U132 ( .A0(N73), .A1(n9), .B0(N40), .B1(n69), .Y(n275) );
  NAND4X1 U133 ( .A(n226), .B(n227), .C(n228), .D(n229), .Y(alu_result[19]) );
  AOI22X1 U134 ( .A0(n46), .A1(n230), .B0(source2[19]), .B1(n231), .Y(n229) );
  AOI22X1 U135 ( .A0(rotate_tmp[19]), .A1(n85), .B0(N208), .B1(n10), .Y(n227)
         );
  AOI22X1 U136 ( .A0(N80), .A1(n9), .B0(N47), .B1(n69), .Y(n226) );
  NAND4X1 U137 ( .A(n212), .B(n213), .C(n214), .D(n215), .Y(alu_result[20]) );
  AOI22X1 U138 ( .A0(n47), .A1(n216), .B0(source2[20]), .B1(n217), .Y(n215) );
  AOI22X1 U139 ( .A0(rotate_tmp[20]), .A1(n85), .B0(N209), .B1(n10), .Y(n213)
         );
  AOI22X1 U140 ( .A0(N81), .A1(n9), .B0(N48), .B1(n69), .Y(n212) );
  NAND4X1 U141 ( .A(n268), .B(n269), .C(n270), .D(n271), .Y(alu_result[13]) );
  AOI22X1 U142 ( .A0(n40), .A1(n272), .B0(source2[13]), .B1(n273), .Y(n271) );
  AOI22X1 U143 ( .A0(rotate_tmp[13]), .A1(n85), .B0(N202), .B1(n10), .Y(n269)
         );
  AOI22X1 U144 ( .A0(N74), .A1(n9), .B0(N41), .B1(n69), .Y(n268) );
  NAND4X1 U145 ( .A(n240), .B(n241), .C(n242), .D(n243), .Y(alu_result[17]) );
  AOI22X1 U146 ( .A0(n44), .A1(n244), .B0(source2[17]), .B1(n245), .Y(n243) );
  AOI22X1 U147 ( .A0(rotate_tmp[17]), .A1(n85), .B0(N206), .B1(n10), .Y(n241)
         );
  AOI22X1 U148 ( .A0(N78), .A1(n9), .B0(N45), .B1(n69), .Y(n240) );
  NAND4X1 U149 ( .A(n282), .B(n283), .C(n284), .D(n285), .Y(alu_result[11]) );
  AOI22X1 U150 ( .A0(n38), .A1(n286), .B0(source2[11]), .B1(n287), .Y(n285) );
  AOI22X1 U151 ( .A0(rotate_tmp[11]), .A1(n85), .B0(N200), .B1(n10), .Y(n283)
         );
  AOI22X1 U152 ( .A0(N72), .A1(n9), .B0(N39), .B1(n69), .Y(n282) );
  NAND4X1 U153 ( .A(n254), .B(n255), .C(n256), .D(n257), .Y(alu_result[15]) );
  AOI22X1 U154 ( .A0(n42), .A1(n258), .B0(source2[15]), .B1(n259), .Y(n257) );
  AOI22X1 U155 ( .A0(rotate_tmp[15]), .A1(n85), .B0(N204), .B1(n10), .Y(n255)
         );
  AOI22X1 U156 ( .A0(N76), .A1(n9), .B0(N43), .B1(n69), .Y(n254) );
  NAND4X1 U157 ( .A(n261), .B(n262), .C(n263), .D(n264), .Y(alu_result[14]) );
  AOI22X1 U158 ( .A0(n41), .A1(n265), .B0(source2[14]), .B1(n266), .Y(n264) );
  AOI22X1 U159 ( .A0(rotate_tmp[14]), .A1(n85), .B0(N203), .B1(n10), .Y(n262)
         );
  AOI22X1 U160 ( .A0(N75), .A1(n9), .B0(N42), .B1(n69), .Y(n261) );
  NAND4X1 U161 ( .A(n296), .B(n297), .C(n298), .D(n299), .Y(alu_result[0]) );
  AOI22X1 U162 ( .A0(n27), .A1(n300), .B0(n14), .B1(n301), .Y(n299) );
  AOI22X1 U163 ( .A0(N61), .A1(n9), .B0(N28), .B1(n69), .Y(n296) );
  AOI22X1 U164 ( .A0(rotate_tmp[0]), .A1(n85), .B0(N189), .B1(n10), .Y(n297)
         );
  NAND4X1 U165 ( .A(n219), .B(n220), .C(n221), .D(n222), .Y(alu_result[1]) );
  AOI22X1 U166 ( .A0(n28), .A1(n223), .B0(n15), .B1(n224), .Y(n222) );
  AOI22X1 U167 ( .A0(N62), .A1(n9), .B0(N29), .B1(n69), .Y(n219) );
  AOI22X1 U168 ( .A0(rotate_tmp[1]), .A1(n85), .B0(N190), .B1(n10), .Y(n220)
         );
  NAND4X1 U169 ( .A(n142), .B(n143), .C(n144), .D(n145), .Y(alu_result[2]) );
  AOI22X1 U170 ( .A0(n29), .A1(n146), .B0(n21), .B1(n147), .Y(n145) );
  AOI22X1 U171 ( .A0(N63), .A1(n9), .B0(N30), .B1(n69), .Y(n142) );
  AOI22X1 U172 ( .A0(rotate_tmp[2]), .A1(n85), .B0(N191), .B1(n10), .Y(n143)
         );
  NAND4X1 U173 ( .A(n122), .B(n123), .C(n124), .D(n125), .Y(alu_result[3]) );
  AOI22X1 U174 ( .A0(n30), .A1(n126), .B0(n23), .B1(n127), .Y(n125) );
  AOI22X1 U175 ( .A0(N64), .A1(n9), .B0(N31), .B1(n69), .Y(n122) );
  AOI22X1 U176 ( .A0(rotate_tmp[3]), .A1(n85), .B0(N192), .B1(n10), .Y(n123)
         );
  NAND4X1 U177 ( .A(n115), .B(n116), .C(n117), .D(n118), .Y(alu_result[4]) );
  AOI22X1 U178 ( .A0(n31), .A1(n119), .B0(n24), .B1(n120), .Y(n118) );
  AOI22X1 U179 ( .A0(N65), .A1(n9), .B0(N32), .B1(n69), .Y(n115) );
  AOI22X1 U180 ( .A0(rotate_tmp[4]), .A1(n85), .B0(N193), .B1(n10), .Y(n116)
         );
  NAND4X1 U181 ( .A(n108), .B(n109), .C(n110), .D(n111), .Y(alu_result[5]) );
  AOI22X1 U182 ( .A0(n32), .A1(n112), .B0(n25), .B1(n113), .Y(n111) );
  AOI22X1 U183 ( .A0(N66), .A1(n9), .B0(N33), .B1(n69), .Y(n108) );
  AOI22X1 U184 ( .A0(rotate_tmp[5]), .A1(n85), .B0(N194), .B1(n10), .Y(n109)
         );
  AOI22X1 U185 ( .A0(N253), .A1(n5), .B0(N221), .B1(n84), .Y(n298) );
  NAND2BX1 U186 ( .AN(n24), .B(n358), .Y(n423) );
  NAND2BX1 U187 ( .AN(n24), .B(n357), .Y(n422) );
  NAND2X1 U188 ( .A(n357), .B(n24), .Y(n433) );
  OR2X2 U189 ( .A(n204), .B(n24), .Y(n431) );
  OAI221XL U190 ( .A0(n33), .A1(n2), .B0(n11), .B1(n342), .C0(n6), .Y(n106) );
  OAI221XL U191 ( .A0(n34), .A1(n2), .B0(n11), .B1(n341), .C0(n6), .Y(n99) );
  OAI221XL U192 ( .A0(n35), .A1(n2), .B0(n11), .B1(n315), .C0(n6), .Y(n92) );
  OAI221XL U193 ( .A0(n36), .A1(n2), .B0(n314), .B1(n11), .C0(n6), .Y(n77) );
  OAI221XL U194 ( .A0(n37), .A1(n2), .B0(n11), .B1(n339), .C0(n6), .Y(n294) );
  OAI221XL U195 ( .A0(n38), .A1(n2), .B0(n11), .B1(n338), .C0(n6), .Y(n287) );
  OAI221XL U196 ( .A0(n39), .A1(n2), .B0(n11), .B1(n281), .C0(n6), .Y(n280) );
  OAI221XL U197 ( .A0(n40), .A1(n2), .B0(n11), .B1(n274), .C0(n6), .Y(n273) );
  OAI221XL U198 ( .A0(n41), .A1(n2), .B0(n11), .B1(n328), .C0(n6), .Y(n266) );
  OAI221XL U199 ( .A0(n42), .A1(n2), .B0(n11), .B1(n327), .C0(n6), .Y(n259) );
  OAI221XL U200 ( .A0(n43), .A1(n2), .B0(n11), .B1(n260), .C0(n6), .Y(n252) );
  OAI221XL U201 ( .A0(n44), .A1(n2), .B0(n11), .B1(n253), .C0(n6), .Y(n245) );
  OAI221XL U202 ( .A0(n45), .A1(n2), .B0(n11), .B1(n325), .C0(n6), .Y(n238) );
  OAI221XL U203 ( .A0(n46), .A1(n2), .B0(n11), .B1(n451), .C0(n6), .Y(n231) );
  OAI221XL U204 ( .A0(n47), .A1(n2), .B0(n11), .B1(n446), .C0(n6), .Y(n217) );
  OAI221XL U205 ( .A0(n48), .A1(n2), .B0(n11), .B1(n445), .C0(n6), .Y(n210) );
  OAI221XL U206 ( .A0(n49), .A1(n2), .B0(n11), .B1(n457), .C0(n6), .Y(n203) );
  OAI221XL U207 ( .A0(n50), .A1(n2), .B0(n11), .B1(n456), .C0(n6), .Y(n196) );
  OAI221XL U208 ( .A0(n51), .A1(n2), .B0(n11), .B1(n443), .C0(n6), .Y(n189) );
  OAI221XL U209 ( .A0(n52), .A1(n2), .B0(n11), .B1(n442), .C0(n6), .Y(n182) );
  OAI221XL U210 ( .A0(n53), .A1(n2), .B0(n11), .B1(n454), .C0(n6), .Y(n175) );
  OAI221XL U211 ( .A0(n54), .A1(n2), .B0(n11), .B1(n453), .C0(n6), .Y(n168) );
  OAI221XL U212 ( .A0(n55), .A1(n2), .B0(n11), .B1(n449), .C0(n6), .Y(n161) );
  OAI221XL U213 ( .A0(n56), .A1(n2), .B0(n11), .B1(n448), .C0(n6), .Y(n154) );
  OAI221XL U214 ( .A0(n57), .A1(n2), .B0(n11), .B1(n435), .C0(n6), .Y(n140) );
  OAI221XL U215 ( .A0(n58), .A1(n2), .B0(n70), .B1(n11), .C0(n6), .Y(n134) );
  NAND2X1 U216 ( .A(n303), .B(n310), .Y(n307) );
  OAI21XL U217 ( .A0(source2[9]), .A1(n2), .B0(n62), .Y(n76) );
  OAI21XL U218 ( .A0(source2[8]), .A1(n2), .B0(n62), .Y(n91) );
  OAI21XL U219 ( .A0(source2[7]), .A1(n2), .B0(n62), .Y(n98) );
  OAI21XL U220 ( .A0(source2[28]), .A1(n2), .B0(n62), .Y(n160) );
  OAI21XL U221 ( .A0(source2[27]), .A1(n2), .B0(n62), .Y(n167) );
  OAI21XL U222 ( .A0(source2[26]), .A1(n2), .B0(n62), .Y(n174) );
  OAI21XL U223 ( .A0(source2[22]), .A1(n2), .B0(n62), .Y(n202) );
  NAND2X1 U224 ( .A(n309), .B(n311), .Y(n306) );
  OAI21XL U225 ( .A0(source2[25]), .A1(n2), .B0(n62), .Y(n181) );
  OAI21XL U226 ( .A0(source2[29]), .A1(n2), .B0(n62), .Y(n153) );
  OAI21XL U227 ( .A0(source2[6]), .A1(n2), .B0(n62), .Y(n105) );
  OAI21XL U228 ( .A0(source2[30]), .A1(n2), .B0(n62), .Y(n139) );
  OAI21XL U229 ( .A0(source2[24]), .A1(n2), .B0(n62), .Y(n188) );
  OAI21XL U230 ( .A0(source2[23]), .A1(n2), .B0(n62), .Y(n195) );
  OAI21XL U231 ( .A0(source2[10]), .A1(n2), .B0(n62), .Y(n293) );
  OAI21XL U232 ( .A0(source2[18]), .A1(n2), .B0(n62), .Y(n237) );
  OAI21XL U233 ( .A0(source2[16]), .A1(n2), .B0(n62), .Y(n251) );
  OAI21XL U234 ( .A0(source2[21]), .A1(n2), .B0(n62), .Y(n209) );
  OAI21XL U235 ( .A0(source2[12]), .A1(n2), .B0(n62), .Y(n279) );
  OAI21XL U236 ( .A0(source2[19]), .A1(n2), .B0(n62), .Y(n230) );
  OAI21XL U237 ( .A0(source2[20]), .A1(n2), .B0(n62), .Y(n216) );
  OAI21XL U238 ( .A0(source2[13]), .A1(n2), .B0(n62), .Y(n272) );
  OAI21XL U239 ( .A0(source2[17]), .A1(n2), .B0(n62), .Y(n244) );
  OAI21XL U240 ( .A0(source2[11]), .A1(n2), .B0(n62), .Y(n286) );
  OAI21XL U241 ( .A0(source2[15]), .A1(n2), .B0(n62), .Y(n258) );
  OAI21XL U242 ( .A0(source2[14]), .A1(n2), .B0(n62), .Y(n265) );
  OAI21XL U243 ( .A0(n14), .A1(n2), .B0(n62), .Y(n300) );
  OAI21XL U244 ( .A0(n15), .A1(n2), .B0(n62), .Y(n223) );
  OAI21XL U245 ( .A0(n21), .A1(n2), .B0(n62), .Y(n146) );
  OAI21XL U246 ( .A0(n25), .A1(n2), .B0(n62), .Y(n112) );
  OAI21XL U247 ( .A0(n26), .A1(n2), .B0(n62), .Y(n133) );
  OAI21XL U248 ( .A0(n23), .A1(n2), .B0(n62), .Y(n126) );
  OAI21XL U249 ( .A0(n24), .A1(n2), .B0(n62), .Y(n119) );
  NOR2BX1 U250 ( .AN(n304), .B(n307), .Y(n69) );
  OAI221XL U251 ( .A0(n306), .A1(n307), .B0(n308), .B1(n309), .C0(n6), .Y(n305) );
  INVX1 U252 ( .A(n307), .Y(n308) );
  INVX1 U253 ( .A(n58), .Y(n70) );
  OAI221XL U254 ( .A0(n30), .A1(n2), .B0(n11), .B1(n333), .C0(n6), .Y(n127) );
  OAI221XL U255 ( .A0(n31), .A1(n2), .B0(n11), .B1(n318), .C0(n6), .Y(n120) );
  OAI221XL U256 ( .A0(n32), .A1(n2), .B0(n11), .B1(n317), .C0(n6), .Y(n113) );
  OAI221XL U257 ( .A0(n29), .A1(n2), .B0(n11), .B1(n334), .C0(n6), .Y(n147) );
  OAI221XL U258 ( .A0(n28), .A1(n2), .B0(n11), .B1(n211), .C0(n6), .Y(n224) );
  OAI221XL U259 ( .A0(n27), .A1(n2), .B0(n11), .B1(n335), .C0(n6), .Y(n301) );
  AOI33X1 U260 ( .A0(n9), .A1(n70), .A2(N285), .B0(n58), .B1(n71), .B2(n69), 
        .Y(n64) );
  INVX1 U261 ( .A(N59), .Y(n71) );
  AOI33X1 U262 ( .A0(n9), .A1(n68), .A2(n58), .B0(n69), .B1(n70), .B2(N59), 
        .Y(n66) );
  INVX1 U263 ( .A(N285), .Y(n68) );
  OAI22X1 U264 ( .A0(n64), .A1(n65), .B0(n26), .B1(n66), .Y(over_flow) );
  INVX1 U265 ( .A(n26), .Y(n65) );
  AND2X2 U266 ( .A(sv[0]), .B(ls_w_mode), .Y(N14) );
  NAND2BX1 U267 ( .AN(sv[1]), .B(ls_w_mode), .Y(N15) );
  BUFX3 U268 ( .A(source2[4]), .Y(n24) );
  BUFX3 U269 ( .A(source2[2]), .Y(n21) );
  BUFX3 U270 ( .A(source2[3]), .Y(n23) );
  BUFX3 U271 ( .A(source1[3]), .Y(n30) );
  BUFX3 U272 ( .A(source1[4]), .Y(n31) );
  BUFX3 U273 ( .A(source1[5]), .Y(n32) );
  BUFX3 U274 ( .A(source1[6]), .Y(n33) );
  BUFX3 U275 ( .A(source1[7]), .Y(n34) );
  BUFX3 U276 ( .A(source1[8]), .Y(n35) );
  BUFX3 U277 ( .A(source1[9]), .Y(n36) );
  BUFX3 U278 ( .A(source1[2]), .Y(n29) );
  BUFX3 U279 ( .A(source1[1]), .Y(n28) );
  BUFX3 U280 ( .A(source2[1]), .Y(n15) );
  BUFX3 U281 ( .A(source1[0]), .Y(n27) );
  BUFX3 U282 ( .A(source2[5]), .Y(n25) );
  BUFX3 U283 ( .A(source2[0]), .Y(n14) );
  BUFX3 U284 ( .A(source1[14]), .Y(n41) );
  BUFX3 U285 ( .A(source2[31]), .Y(n26) );
  BUFX3 U286 ( .A(source1[15]), .Y(n42) );
  BUFX3 U287 ( .A(source1[16]), .Y(n43) );
  BUFX3 U288 ( .A(source1[10]), .Y(n37) );
  BUFX3 U289 ( .A(source1[11]), .Y(n38) );
  BUFX3 U290 ( .A(source1[12]), .Y(n39) );
  BUFX3 U291 ( .A(source1[13]), .Y(n40) );
  BUFX3 U292 ( .A(source1[17]), .Y(n44) );
  BUFX3 U293 ( .A(source1[18]), .Y(n45) );
  BUFX3 U294 ( .A(source1[19]), .Y(n46) );
  BUFX3 U295 ( .A(source1[20]), .Y(n47) );
  BUFX3 U296 ( .A(source1[29]), .Y(n56) );
  BUFX3 U297 ( .A(source1[31]), .Y(n58) );
  BUFX3 U298 ( .A(source1[30]), .Y(n57) );
  BUFX3 U299 ( .A(source1[22]), .Y(n49) );
  BUFX3 U300 ( .A(source1[23]), .Y(n50) );
  BUFX3 U301 ( .A(source1[24]), .Y(n51) );
  BUFX3 U302 ( .A(source1[21]), .Y(n48) );
  BUFX3 U303 ( .A(source1[25]), .Y(n52) );
  BUFX3 U304 ( .A(source1[26]), .Y(n53) );
  BUFX3 U305 ( .A(source1[27]), .Y(n54) );
  BUFX3 U306 ( .A(source1[28]), .Y(n55) );
  NOR2X1 U307 ( .A(n311), .B(funct[3]), .Y(n304) );
  NOR3X1 U308 ( .A(n307), .B(funct[0]), .C(n309), .Y(n85) );
  INVX1 U309 ( .A(funct[1]), .Y(n310) );
  INVX1 U310 ( .A(funct[2]), .Y(n303) );
  INVX1 U311 ( .A(funct[3]), .Y(n309) );
  INVX1 U312 ( .A(funct[0]), .Y(n311) );
  AND3X2 U313 ( .A(n304), .B(funct[1]), .C(funct[2]), .Y(n84) );
  NOR3X1 U314 ( .A(source2[13]), .B(source2[15]), .C(source2[14]), .Y(n63) );
  NOR4BX1 U315 ( .AN(n63), .B(source2[12]), .C(source2[10]), .D(source2[11]), 
        .Y(n83) );
  NOR4X1 U316 ( .A(source2[22]), .B(source2[21]), .C(source2[20]), .D(
        source2[19]), .Y(n67) );
  NOR4BX1 U317 ( .AN(n67), .B(source2[18]), .C(source2[16]), .D(source2[17]), 
        .Y(n82) );
  NOR3X1 U318 ( .A(source2[26]), .B(source2[28]), .C(source2[27]), .Y(n78) );
  NOR4BX1 U319 ( .AN(n78), .B(source2[25]), .C(source2[23]), .D(source2[24]), 
        .Y(n81) );
  NOR4X1 U320 ( .A(source2[9]), .B(source2[8]), .C(source2[7]), .D(source2[6]), 
        .Y(n79) );
  NOR4BX1 U321 ( .AN(n79), .B(n26), .C(source2[29]), .D(source2[30]), .Y(n80)
         );
  NAND4X1 U322 ( .A(n83), .B(n82), .C(n81), .D(n80), .Y(n356) );
  NOR2X1 U323 ( .A(n356), .B(n25), .Y(n358) );
  NOR2BX1 U324 ( .AN(n25), .B(n356), .Y(n357) );
  NOR2X1 U325 ( .A(n358), .B(n357), .Y(n204) );
  INVX1 U326 ( .A(n14), .Y(n86) );
  NOR2X1 U327 ( .A(n86), .B(n15), .Y(n331) );
  INVX1 U328 ( .A(n32), .Y(n317) );
  INVX1 U329 ( .A(n33), .Y(n342) );
  NAND2X1 U330 ( .A(n15), .B(n14), .Y(n336) );
  AOI22X1 U331 ( .A0(n34), .A1(n59), .B0(n31), .B1(n1), .Y(n93) );
  OAI221XL U332 ( .A0(n61), .A1(n317), .B0(n60), .B1(n342), .C0(n93), .Y(n393)
         );
  INVX1 U333 ( .A(n21), .Y(n107) );
  INVX1 U334 ( .A(n28), .Y(n211) );
  INVX1 U335 ( .A(n29), .Y(n334) );
  AOI22X1 U336 ( .A0(n30), .A1(n59), .B0(n27), .B1(n1), .Y(n100) );
  OAI221XL U337 ( .A0(n61), .A1(n211), .B0(n60), .B1(n334), .C0(n100), .Y(n392) );
  INVX1 U338 ( .A(n23), .Y(n302) );
  INVX1 U339 ( .A(n40), .Y(n274) );
  INVX1 U340 ( .A(n41), .Y(n328) );
  AOI22X1 U341 ( .A0(n42), .A1(n59), .B0(n39), .B1(n1), .Y(n114) );
  OAI221XL U342 ( .A0(n61), .A1(n274), .B0(n60), .B1(n328), .C0(n114), .Y(n399) );
  INVX1 U343 ( .A(n36), .Y(n314) );
  INVX1 U344 ( .A(n37), .Y(n339) );
  AOI22X1 U345 ( .A0(n38), .A1(n59), .B0(n35), .B1(n1), .Y(n121) );
  OAI221XL U346 ( .A0(n61), .A1(n314), .B0(n60), .B1(n339), .C0(n121), .Y(n398) );
  AOI22X1 U347 ( .A0(n4), .A1(n399), .B0(n8), .B1(n398), .Y(n128) );
  INVX1 U348 ( .A(n128), .Y(n141) );
  AOI221X1 U349 ( .A0(n393), .A1(n7), .B0(n392), .B1(n3), .C0(n141), .Y(n354)
         );
  INVX1 U350 ( .A(n44), .Y(n253) );
  AOI22X1 U351 ( .A0(n46), .A1(n59), .B0(n43), .B1(n1), .Y(n148) );
  OAI221XL U352 ( .A0(n61), .A1(n253), .B0(n60), .B1(n325), .C0(n148), .Y(n394) );
  AOI22X1 U353 ( .A0(n7), .A1(n395), .B0(n3), .B1(n394), .Y(n155) );
  INVX1 U354 ( .A(n155), .Y(n162) );
  AOI221X1 U355 ( .A0(n390), .A1(n4), .B0(n391), .B1(n8), .C0(n162), .Y(n355)
         );
  MX2X1 U356 ( .A(n354), .B(n355), .S0(n24), .Y(n169) );
  NOR2X1 U357 ( .A(n204), .B(n169), .Y(rotate_tmp[0]) );
  INVX1 U358 ( .A(n42), .Y(n327) );
  INVX1 U359 ( .A(n43), .Y(n260) );
  AOI22X1 U360 ( .A0(n44), .A1(n59), .B0(n41), .B1(n1), .Y(n176) );
  OAI221XL U361 ( .A0(n61), .A1(n327), .B0(n60), .B1(n260), .C0(n176), .Y(n375) );
  INVX1 U362 ( .A(n38), .Y(n338) );
  INVX1 U363 ( .A(n39), .Y(n281) );
  AOI22X1 U364 ( .A0(n40), .A1(n59), .B0(n37), .B1(n1), .Y(n183) );
  OAI221XL U365 ( .A0(n61), .A1(n338), .B0(n60), .B1(n281), .C0(n183), .Y(n380) );
  AOI22X1 U366 ( .A0(n4), .A1(n373), .B0(n8), .B1(n376), .Y(n190) );
  INVX1 U367 ( .A(n190), .Y(n197) );
  AOI221X1 U368 ( .A0(n375), .A1(n7), .B0(n380), .B1(n3), .C0(n197), .Y(n411)
         );
  INVX1 U369 ( .A(n27), .Y(n335) );
  INVX1 U370 ( .A(n34), .Y(n341) );
  INVX1 U371 ( .A(n35), .Y(n315) );
  AOI22X1 U372 ( .A0(n36), .A1(n59), .B0(n33), .B1(n1), .Y(n218) );
  OAI221XL U373 ( .A0(n61), .A1(n341), .B0(n60), .B1(n315), .C0(n218), .Y(n379) );
  INVX1 U374 ( .A(n30), .Y(n333) );
  INVX1 U375 ( .A(n31), .Y(n318) );
  AOI22X1 U376 ( .A0(n32), .A1(n59), .B0(n29), .B1(n1), .Y(n225) );
  OAI221XL U377 ( .A0(n61), .A1(n333), .B0(n60), .B1(n318), .C0(n225), .Y(n374) );
  AOI22X1 U378 ( .A0(n4), .A1(n379), .B0(n8), .B1(n374), .Y(n232) );
  INVX1 U379 ( .A(n232), .Y(n239) );
  AOI22X1 U380 ( .A0(n45), .A1(n59), .B0(n42), .B1(n1), .Y(n246) );
  OAI221XL U381 ( .A0(n61), .A1(n260), .B0(n60), .B1(n253), .C0(n246), .Y(n384) );
  AOI22X1 U382 ( .A0(n41), .A1(n59), .B0(n38), .B1(n1), .Y(n267) );
  OAI221XL U383 ( .A0(n61), .A1(n281), .B0(n60), .B1(n274), .C0(n267), .Y(n389) );
  AOI22X1 U384 ( .A0(n4), .A1(n382), .B0(n8), .B1(n385), .Y(n288) );
  INVX1 U385 ( .A(n288), .Y(n295) );
  AOI221X1 U386 ( .A0(n384), .A1(n7), .B0(n389), .B1(n3), .C0(n295), .Y(n412)
         );
  AOI22X1 U387 ( .A0(n28), .A1(n12), .B0(n29), .B1(n59), .Y(n312) );
  AOI22X1 U388 ( .A0(n37), .A1(n59), .B0(n34), .B1(n1), .Y(n313) );
  OAI221XL U389 ( .A0(n61), .A1(n315), .B0(n60), .B1(n314), .C0(n313), .Y(n388) );
  AOI22X1 U390 ( .A0(n33), .A1(n59), .B0(n30), .B1(n1), .Y(n316) );
  OAI221XL U391 ( .A0(n61), .A1(n318), .B0(n60), .B1(n317), .C0(n316), .Y(n383) );
  AOI22X1 U392 ( .A0(n4), .A1(n388), .B0(n8), .B1(n383), .Y(n319) );
  INVX1 U393 ( .A(n319), .Y(n320) );
  AOI22X1 U394 ( .A0(n4), .A1(n391), .B0(n8), .B1(n395), .Y(n321) );
  INVX1 U395 ( .A(n321), .Y(n322) );
  AOI221X1 U396 ( .A0(n394), .A1(n7), .B0(n399), .B1(n3), .C0(n322), .Y(n413)
         );
  NAND2BX1 U397 ( .AN(n433), .B(n3), .Y(n353) );
  AOI22X1 U398 ( .A0(n4), .A1(n398), .B0(n8), .B1(n393), .Y(n323) );
  INVX1 U399 ( .A(n323), .Y(n324) );
  AOI22X1 U400 ( .A0(n43), .A1(n59), .B0(n40), .B1(n1), .Y(n326) );
  OAI221XL U401 ( .A0(n61), .A1(n328), .B0(n60), .B1(n327), .C0(n326), .Y(n410) );
  AOI22X1 U402 ( .A0(n4), .A1(n404), .B0(n8), .B1(n406), .Y(n329) );
  INVX1 U403 ( .A(n329), .Y(n330) );
  AOI221X1 U404 ( .A0(n405), .A1(n7), .B0(n410), .B1(n3), .C0(n330), .Y(n414)
         );
  AOI22X1 U405 ( .A0(n31), .A1(n59), .B0(n28), .B1(n1), .Y(n332) );
  OAI221XL U406 ( .A0(n61), .A1(n334), .B0(n60), .B1(n333), .C0(n332), .Y(n400) );
  AOI22X1 U407 ( .A0(n39), .A1(n59), .B0(n36), .B1(n1), .Y(n337) );
  OAI221XL U408 ( .A0(n61), .A1(n339), .B0(n60), .B1(n338), .C0(n337), .Y(n409) );
  AOI22X1 U409 ( .A0(n35), .A1(n59), .B0(n32), .B1(n1), .Y(n340) );
  OAI221XL U410 ( .A0(n61), .A1(n342), .B0(n60), .B1(n341), .C0(n340), .Y(n401) );
  AOI22X1 U411 ( .A0(n4), .A1(n409), .B0(n8), .B1(n401), .Y(n343) );
  INVX1 U412 ( .A(n343), .Y(n344) );
  AOI22X1 U413 ( .A0(n7), .A1(n376), .B0(n3), .B1(n375), .Y(n345) );
  INVX1 U414 ( .A(n345), .Y(n346) );
  AOI221X1 U415 ( .A0(n372), .A1(n4), .B0(n373), .B1(n8), .C0(n346), .Y(n418)
         );
  AOI22X1 U416 ( .A0(n4), .A1(n380), .B0(n8), .B1(n379), .Y(n347) );
  INVX1 U417 ( .A(n347), .Y(n348) );
  AOI22X1 U418 ( .A0(n7), .A1(n385), .B0(n3), .B1(n384), .Y(n349) );
  INVX1 U419 ( .A(n349), .Y(n350) );
  AOI221X1 U420 ( .A0(n381), .A1(n4), .B0(n382), .B1(n8), .C0(n350), .Y(n419)
         );
  AOI22X1 U421 ( .A0(n4), .A1(n389), .B0(n8), .B1(n388), .Y(n351) );
  INVX1 U422 ( .A(n351), .Y(n352) );
  OAI32X1 U423 ( .A0(n356), .A1(n24), .A2(n355), .B0(n354), .B1(n13), .Y(
        rotate_tmp[16]) );
  AOI22X1 U424 ( .A0(n4), .A1(n410), .B0(n8), .B1(n409), .Y(n359) );
  INVX1 U425 ( .A(n359), .Y(n360) );
  AOI221X1 U426 ( .A0(n401), .A1(n7), .B0(n400), .B1(n3), .C0(n360), .Y(n365)
         );
  AOI22X1 U427 ( .A0(n4), .A1(n375), .B0(n8), .B1(n380), .Y(n361) );
  INVX1 U428 ( .A(n361), .Y(n362) );
  AOI221X1 U429 ( .A0(n379), .A1(n7), .B0(n374), .B1(n3), .C0(n362), .Y(n415)
         );
  AOI22X1 U430 ( .A0(n4), .A1(n384), .B0(n8), .B1(n389), .Y(n363) );
  INVX1 U431 ( .A(n363), .Y(n364) );
  AOI221X1 U432 ( .A0(n388), .A1(n7), .B0(n383), .B1(n3), .C0(n364), .Y(n421)
         );
  AOI21X1 U433 ( .A0(n423), .A1(n422), .B0(n365), .Y(n366) );
  INVX1 U434 ( .A(n366), .Y(n367) );
  AOI22X1 U435 ( .A0(n4), .A1(n394), .B0(n8), .B1(n399), .Y(n368) );
  INVX1 U436 ( .A(n368), .Y(n369) );
  AOI221X1 U437 ( .A0(n398), .A1(n7), .B0(n393), .B1(n3), .C0(n369), .Y(n426)
         );
  AOI22X1 U438 ( .A0(n4), .A1(n405), .B0(n8), .B1(n410), .Y(n370) );
  INVX1 U439 ( .A(n370), .Y(n371) );
  AOI221X1 U440 ( .A0(n409), .A1(n7), .B0(n401), .B1(n3), .C0(n371), .Y(n427)
         );
  AOI22X1 U441 ( .A0(n4), .A1(n376), .B0(n8), .B1(n375), .Y(n377) );
  INVX1 U442 ( .A(n377), .Y(n378) );
  AOI221X1 U443 ( .A0(n380), .A1(n7), .B0(n379), .B1(n3), .C0(n378), .Y(n428)
         );
  AOI22X1 U444 ( .A0(n4), .A1(n385), .B0(n8), .B1(n384), .Y(n386) );
  INVX1 U445 ( .A(n386), .Y(n387) );
  AOI221X1 U446 ( .A0(n389), .A1(n7), .B0(n388), .B1(n3), .C0(n387), .Y(n429)
         );
  AOI22X1 U447 ( .A0(n4), .A1(n395), .B0(n8), .B1(n394), .Y(n396) );
  INVX1 U448 ( .A(n396), .Y(n397) );
  AOI221X1 U449 ( .A0(n399), .A1(n7), .B0(n398), .B1(n3), .C0(n397), .Y(n430)
         );
  AOI22X1 U450 ( .A0(n4), .A1(n401), .B0(n8), .B1(n400), .Y(n402) );
  INVX1 U451 ( .A(n402), .Y(n403) );
  AOI22X1 U452 ( .A0(n4), .A1(n406), .B0(n8), .B1(n405), .Y(n407) );
  INVX1 U453 ( .A(n407), .Y(n408) );
  AOI221X1 U454 ( .A0(n410), .A1(n7), .B0(n409), .B1(n3), .C0(n408), .Y(n432)
         );
  NAND2BX1 U455 ( .AN(n422), .B(n3), .Y(n420) );
  AOI21X1 U456 ( .A0(n423), .A1(n422), .B0(n415), .Y(n416) );
  INVX1 U457 ( .A(n416), .Y(n417) );
  AOI21X1 U458 ( .A0(n423), .A1(n422), .B0(n421), .Y(n424) );
  INVX1 U459 ( .A(n424), .Y(n425) );
  INVX1 U460 ( .A(n45), .Y(n325) );
  INVX1 U461 ( .A(n46), .Y(n451) );
  INVX1 U462 ( .A(n47), .Y(n446) );
  OAI221XL U463 ( .A0(n61), .A1(n325), .B0(n60), .B1(n451), .C0(n450), .Y(n405) );
  AOI22X1 U464 ( .A0(n47), .A1(n59), .B0(n44), .B1(n1), .Y(n450) );
  INVX1 U465 ( .A(n48), .Y(n445) );
  OAI221XL U466 ( .A0(n61), .A1(n451), .B0(n60), .B1(n446), .C0(n440), .Y(n376) );
  AOI22X1 U467 ( .A0(n48), .A1(n59), .B0(n45), .B1(n1), .Y(n440) );
  INVX1 U468 ( .A(n49), .Y(n457) );
  OAI221XL U469 ( .A0(n61), .A1(n446), .B0(n60), .B1(n445), .C0(n444), .Y(n385) );
  AOI22X1 U470 ( .A0(n59), .A1(n49), .B0(n46), .B1(n1), .Y(n444) );
  OAI221XL U471 ( .A0(n61), .A1(n445), .B0(n457), .B1(n60), .C0(n437), .Y(n395) );
  AOI22X1 U472 ( .A0(n59), .A1(n50), .B0(n47), .B1(n1), .Y(n437) );
  INVX1 U473 ( .A(n50), .Y(n456) );
  INVX1 U474 ( .A(n51), .Y(n443) );
  OAI221XL U475 ( .A0(n61), .A1(n457), .B0(n60), .B1(n456), .C0(n455), .Y(n406) );
  AOI22X1 U476 ( .A0(n51), .A1(n59), .B0(n48), .B1(n1), .Y(n455) );
  INVX1 U477 ( .A(n52), .Y(n442) );
  OAI221XL U478 ( .A0(n61), .A1(n456), .B0(n60), .B1(n443), .C0(n439), .Y(n373) );
  AOI22X1 U479 ( .A0(n52), .A1(n59), .B0(n1), .B1(n49), .Y(n439) );
  INVX1 U480 ( .A(n53), .Y(n454) );
  INVX1 U481 ( .A(n462), .Y(n464) );
  AOI22X1 U482 ( .A0(n385), .A1(n3), .B0(n382), .B1(n7), .Y(n462) );
  OAI221XL U483 ( .A0(n61), .A1(n443), .B0(n60), .B1(n442), .C0(n441), .Y(n382) );
  AOI22X1 U484 ( .A0(n53), .A1(n59), .B0(n1), .B1(n50), .Y(n441) );
  OAI221XL U485 ( .A0(n61), .A1(n442), .B0(n60), .B1(n454), .C0(n436), .Y(n391) );
  AOI22X1 U486 ( .A0(n54), .A1(n59), .B0(n1), .B1(n51), .Y(n436) );
  INVX1 U487 ( .A(n54), .Y(n453) );
  INVX1 U488 ( .A(n55), .Y(n449) );
  INVX1 U489 ( .A(n468), .Y(n469) );
  AOI22X1 U490 ( .A0(n406), .A1(n3), .B0(n404), .B1(n7), .Y(n468) );
  INVX1 U491 ( .A(n458), .Y(n459) );
  AOI222X1 U492 ( .A0(n406), .A1(n7), .B0(n404), .B1(n8), .C0(n405), .C1(n3), 
        .Y(n458) );
  OAI221XL U493 ( .A0(n61), .A1(n454), .B0(n60), .B1(n453), .C0(n452), .Y(n404) );
  AOI22X1 U494 ( .A0(n55), .A1(n59), .B0(n52), .B1(n1), .Y(n452) );
  INVX1 U495 ( .A(n56), .Y(n448) );
  INVX1 U496 ( .A(n470), .Y(n472) );
  AOI22X1 U497 ( .A0(n373), .A1(n3), .B0(n372), .B1(n7), .Y(n470) );
  INVX1 U498 ( .A(n460), .Y(n461) );
  AOI222X1 U499 ( .A0(n373), .A1(n7), .B0(n372), .B1(n8), .C0(n376), .C1(n3), 
        .Y(n460) );
  OAI221XL U500 ( .A0(n61), .A1(n453), .B0(n60), .B1(n449), .C0(n438), .Y(n372) );
  AOI22X1 U501 ( .A0(n56), .A1(n59), .B0(n53), .B1(n1), .Y(n438) );
  INVX1 U502 ( .A(n57), .Y(n435) );
  INVX1 U503 ( .A(n474), .Y(n476) );
  AOI22X1 U504 ( .A0(n382), .A1(n3), .B0(n381), .B1(n7), .Y(n474) );
  OAI221XL U505 ( .A0(n61), .A1(n449), .B0(n60), .B1(n448), .C0(n447), .Y(n381) );
  AOI22X1 U506 ( .A0(n57), .A1(n59), .B0(n54), .B1(n1), .Y(n447) );
  OAI222XL U507 ( .A0(n506), .A1(n433), .B0(n430), .B1(n431), .C0(n505), .C1(
        n13), .Y(rotate_tmp[8]) );
  OAI222XL U508 ( .A0(n506), .A1(n422), .B0(n505), .B1(n423), .C0(n430), .C1(
        n13), .Y(rotate_tmp[24]) );
  AOI221X1 U509 ( .A0(n393), .A1(n4), .B0(n392), .B1(n8), .C0(n478), .Y(n505)
         );
  INVX1 U510 ( .A(n506), .Y(n478) );
  AOI22X1 U511 ( .A0(n391), .A1(n3), .B0(n390), .B1(n7), .Y(n506) );
  OAI222XL U512 ( .A0(n498), .A1(n433), .B0(n426), .B1(n431), .C0(n497), .C1(
        n13), .Y(rotate_tmp[4]) );
  OAI222XL U513 ( .A0(n498), .A1(n422), .B0(n497), .B1(n423), .C0(n426), .C1(
        n13), .Y(rotate_tmp[20]) );
  AOI21X1 U514 ( .A0(n392), .A1(n4), .B0(n467), .Y(n497) );
  INVX1 U515 ( .A(n498), .Y(n467) );
  AOI222X1 U516 ( .A0(n391), .A1(n7), .B0(n390), .B1(n8), .C0(n395), .C1(n3), 
        .Y(n498) );
  OAI222XL U517 ( .A0(n486), .A1(n423), .B0(n485), .B1(n420), .C0(n413), .C1(
        n13), .Y(rotate_tmp[28]) );
  OAI222XL U518 ( .A0(n413), .A1(n431), .B0(n485), .B1(n353), .C0(n486), .C1(
        n13), .Y(rotate_tmp[12]) );
  AOI221X1 U519 ( .A0(n392), .A1(n7), .B0(n390), .B1(n3), .C0(n324), .Y(n486)
         );
  INVX1 U520 ( .A(n390), .Y(n485) );
  OAI221XL U521 ( .A0(n61), .A1(n448), .B0(n60), .B1(n435), .C0(n434), .Y(n390) );
  AOI22X1 U522 ( .A0(n58), .A1(n59), .B0(n55), .B1(n1), .Y(n434) );
  OAI222XL U523 ( .A0(n492), .A1(n423), .B0(n491), .B1(n420), .C0(n418), .C1(
        n13), .Y(rotate_tmp[30]) );
  OAI222XL U524 ( .A0(n418), .A1(n431), .B0(n491), .B1(n353), .C0(n492), .C1(
        n13), .Y(rotate_tmp[14]) );
  AOI221X1 U525 ( .A0(n374), .A1(n7), .B0(n473), .B1(n3), .C0(n348), .Y(n492)
         );
  OAI222XL U526 ( .A0(n502), .A1(n433), .B0(n428), .B1(n431), .C0(n501), .C1(
        n13), .Y(rotate_tmp[6]) );
  OAI222XL U527 ( .A0(n502), .A1(n422), .B0(n501), .B1(n423), .C0(n428), .C1(
        n13), .Y(rotate_tmp[22]) );
  AOI221X1 U528 ( .A0(n374), .A1(n4), .B0(n473), .B1(n8), .C0(n472), .Y(n501)
         );
  AOI21X1 U529 ( .A0(n471), .A1(n8), .B0(n472), .Y(n502) );
  OAI221XL U530 ( .A0(n490), .A1(n13), .B0(n489), .B1(n433), .C0(n417), .Y(
        rotate_tmp[2]) );
  OAI222XL U531 ( .A0(n489), .A1(n422), .B0(n490), .B1(n423), .C0(n415), .C1(
        n13), .Y(rotate_tmp[18]) );
  AOI21X1 U532 ( .A0(n473), .A1(n4), .B0(n461), .Y(n490) );
  AOI21X1 U533 ( .A0(n471), .A1(n4), .B0(n461), .Y(n489) );
  OAI222XL U534 ( .A0(n482), .A1(n422), .B0(n481), .B1(n423), .C0(n411), .C1(
        n13), .Y(rotate_tmp[26]) );
  OAI222XL U535 ( .A0(n482), .A1(n433), .B0(n411), .B1(n431), .C0(n481), .C1(
        n13), .Y(rotate_tmp[10]) );
  AOI221X1 U536 ( .A0(n473), .A1(n7), .B0(n372), .B1(n3), .C0(n239), .Y(n481)
         );
  OAI221XL U537 ( .A0(n60), .A1(n335), .B0(n336), .B1(n211), .C0(n491), .Y(
        n473) );
  AOI22X1 U538 ( .A0(n372), .A1(n3), .B0(n471), .B1(n7), .Y(n482) );
  INVX1 U539 ( .A(n491), .Y(n471) );
  AOI22X1 U540 ( .A0(n1), .A1(n57), .B0(n331), .B1(n58), .Y(n491) );
  OAI222XL U541 ( .A0(n494), .A1(n423), .B0(n493), .B1(n420), .C0(n419), .C1(
        n13), .Y(rotate_tmp[31]) );
  OAI222XL U542 ( .A0(n419), .A1(n431), .B0(n493), .B1(n353), .C0(n494), .C1(
        n13), .Y(rotate_tmp[15]) );
  AOI221X1 U543 ( .A0(n383), .A1(n7), .B0(n477), .B1(n3), .C0(n352), .Y(n494)
         );
  OAI222XL U544 ( .A0(n504), .A1(n433), .B0(n429), .B1(n431), .C0(n503), .C1(
        n13), .Y(rotate_tmp[7]) );
  OAI222XL U545 ( .A0(n504), .A1(n422), .B0(n503), .B1(n423), .C0(n429), .C1(
        n13), .Y(rotate_tmp[23]) );
  AOI221X1 U546 ( .A0(n383), .A1(n4), .B0(n477), .B1(n8), .C0(n476), .Y(n503)
         );
  AOI21X1 U547 ( .A0(n8), .A1(n475), .B0(n476), .Y(n504) );
  OAI221XL U548 ( .A0(n496), .A1(n13), .B0(n495), .B1(n433), .C0(n425), .Y(
        rotate_tmp[3]) );
  OAI222XL U549 ( .A0(n495), .A1(n422), .B0(n496), .B1(n423), .C0(n421), .C1(
        n13), .Y(rotate_tmp[19]) );
  AOI221X1 U550 ( .A0(n477), .A1(n4), .B0(n381), .B1(n8), .C0(n464), .Y(n496)
         );
  AOI21X1 U551 ( .A0(n23), .A1(n463), .B0(n464), .Y(n495) );
  OAI222XL U552 ( .A0(n484), .A1(n423), .B0(n422), .B1(n483), .C0(n412), .C1(
        n13), .Y(rotate_tmp[27]) );
  OAI222XL U553 ( .A0(n412), .A1(n431), .B0(n433), .B1(n483), .C0(n484), .C1(
        n13), .Y(rotate_tmp[11]) );
  AOI221X1 U554 ( .A0(n477), .A1(n7), .B0(n381), .B1(n3), .C0(n320), .Y(n484)
         );
  OAI211X1 U555 ( .A0(n61), .A1(n335), .B0(n493), .C0(n312), .Y(n477) );
  NAND2X1 U556 ( .A(n463), .B(n302), .Y(n483) );
  MX2X1 U557 ( .A(n381), .B(n475), .S0(n21), .Y(n463) );
  INVX1 U558 ( .A(n493), .Y(n475) );
  NAND2X1 U559 ( .A(n58), .B(n1), .Y(n493) );
  OAI222XL U560 ( .A0(n488), .A1(n423), .B0(n487), .B1(n420), .C0(n414), .C1(
        n13), .Y(rotate_tmp[29]) );
  OAI222XL U561 ( .A0(n508), .A1(n433), .B0(n432), .B1(n431), .C0(n507), .C1(
        n13), .Y(rotate_tmp[9]) );
  OAI222XL U562 ( .A0(n508), .A1(n422), .B0(n507), .B1(n423), .C0(n432), .C1(
        n13), .Y(rotate_tmp[25]) );
  AOI221X1 U563 ( .A0(n480), .A1(n7), .B0(n404), .B1(n3), .C0(n403), .Y(n507)
         );
  AOI22X1 U564 ( .A0(n404), .A1(n3), .B0(n479), .B1(n7), .Y(n508) );
  OAI222XL U565 ( .A0(n500), .A1(n433), .B0(n427), .B1(n431), .C0(n499), .C1(
        n13), .Y(rotate_tmp[5]) );
  OAI222XL U566 ( .A0(n500), .A1(n422), .B0(n499), .B1(n423), .C0(n427), .C1(
        n13), .Y(rotate_tmp[21]) );
  AOI221X1 U567 ( .A0(n400), .A1(n4), .B0(n480), .B1(n8), .C0(n469), .Y(n499)
         );
  AOI21X1 U568 ( .A0(n479), .A1(n8), .B0(n469), .Y(n500) );
  OAI221XL U569 ( .A0(n466), .A1(n13), .B0(n465), .B1(n433), .C0(n367), .Y(
        rotate_tmp[1]) );
  OAI222XL U570 ( .A0(n465), .A1(n422), .B0(n466), .B1(n423), .C0(n365), .C1(
        n13), .Y(rotate_tmp[17]) );
  AOI21X1 U571 ( .A0(n480), .A1(n4), .B0(n459), .Y(n466) );
  AOI21X1 U572 ( .A0(n479), .A1(n4), .B0(n459), .Y(n465) );
  INVX1 U573 ( .A(n487), .Y(n479) );
  OAI222XL U574 ( .A0(n414), .A1(n431), .B0(n487), .B1(n353), .C0(n488), .C1(
        n13), .Y(rotate_tmp[13]) );
  AOI221X1 U575 ( .A0(n400), .A1(n7), .B0(n480), .B1(n3), .C0(n344), .Y(n488)
         );
  OAI21XL U576 ( .A0(n336), .A1(n335), .B0(n487), .Y(n480) );
  AOI222X1 U577 ( .A0(n12), .A1(n58), .B0(n331), .B1(n57), .C0(n1), .C1(n56), 
        .Y(n487) );
endmodule


module IDEX ( ls_w_mode_out, funct_out, sel_in2_out, ena_data_out, data_rw_out, 
        sel_wb_out, reg_rw_out, read_data1_out, read_data2_out, read_data3_out, 
        ext_out, addr_dst_out, ls_w_mode_in, funct_in, sel_in2_in, ena_data_in, 
        data_rw_in, sel_wb_in, reg_rw_in, read_data1_in, read_data2_in, 
        addr_dst_in, read_data3_in, ext_in, clk, rst, addr1_out, addr1_in, 
        addr2_out, addr2_in, inst_out, inst_in, sel_alu_out, sel_alu_in );
  output [3:0] funct_out;
  output [31:0] read_data1_out;
  output [31:0] read_data2_out;
  output [31:0] read_data3_out;
  output [31:0] ext_out;
  output [4:0] addr_dst_out;
  input [3:0] funct_in;
  input [31:0] read_data1_in;
  input [31:0] read_data2_in;
  input [4:0] addr_dst_in;
  input [31:0] read_data3_in;
  input [31:0] ext_in;
  output [4:0] addr1_out;
  input [4:0] addr1_in;
  output [4:0] addr2_out;
  input [4:0] addr2_in;
  output [31:0] inst_out;
  input [31:0] inst_in;
  input ls_w_mode_in, sel_in2_in, ena_data_in, data_rw_in, sel_wb_in,
         reg_rw_in, clk, rst, sel_alu_in;
  output ls_w_mode_out, sel_in2_out, ena_data_out, data_rw_out, sel_wb_out,
         reg_rw_out, sel_alu_out;


  DFFRHQX1 sel_alu_out_reg ( .D(sel_alu_in), .CK(clk), .RN(rst), .Q(
        sel_alu_out) );
  DFFRHQX1 ena_data_out_reg ( .D(ena_data_in), .CK(clk), .RN(rst), .Q(
        ena_data_out) );
  DFFRHQX1 \read_data1_out_reg[31]  ( .D(read_data1_in[31]), .CK(clk), .RN(rst), .Q(read_data1_out[31]) );
  DFFRHQX1 \read_data1_out_reg[30]  ( .D(read_data1_in[30]), .CK(clk), .RN(rst), .Q(read_data1_out[30]) );
  DFFRHQX1 \read_data1_out_reg[29]  ( .D(read_data1_in[29]), .CK(clk), .RN(rst), .Q(read_data1_out[29]) );
  DFFRHQX1 \read_data1_out_reg[28]  ( .D(read_data1_in[28]), .CK(clk), .RN(rst), .Q(read_data1_out[28]) );
  DFFRHQX1 \read_data1_out_reg[27]  ( .D(read_data1_in[27]), .CK(clk), .RN(rst), .Q(read_data1_out[27]) );
  DFFRHQX1 \read_data1_out_reg[26]  ( .D(read_data1_in[26]), .CK(clk), .RN(rst), .Q(read_data1_out[26]) );
  DFFRHQX1 \read_data1_out_reg[25]  ( .D(read_data1_in[25]), .CK(clk), .RN(rst), .Q(read_data1_out[25]) );
  DFFRHQX1 \read_data1_out_reg[24]  ( .D(read_data1_in[24]), .CK(clk), .RN(rst), .Q(read_data1_out[24]) );
  DFFRHQX1 \read_data1_out_reg[23]  ( .D(read_data1_in[23]), .CK(clk), .RN(rst), .Q(read_data1_out[23]) );
  DFFRHQX1 \read_data1_out_reg[22]  ( .D(read_data1_in[22]), .CK(clk), .RN(rst), .Q(read_data1_out[22]) );
  DFFRHQX1 \addr_dst_out_reg[4]  ( .D(addr_dst_in[4]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[4]) );
  DFFRHQX1 \addr_dst_out_reg[2]  ( .D(addr_dst_in[2]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[2]) );
  DFFRHQX1 \addr_dst_out_reg[3]  ( .D(addr_dst_in[3]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[3]) );
  DFFRHQX1 \addr_dst_out_reg[1]  ( .D(addr_dst_in[1]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[1]) );
  DFFRHQX1 \addr_dst_out_reg[0]  ( .D(addr_dst_in[0]), .CK(clk), .RN(rst), .Q(
        addr_dst_out[0]) );
  DFFRHQX1 \funct_out_reg[0]  ( .D(funct_in[0]), .CK(clk), .RN(rst), .Q(
        funct_out[0]) );
  DFFRHQX1 \funct_out_reg[3]  ( .D(funct_in[3]), .CK(clk), .RN(rst), .Q(
        funct_out[3]) );
  DFFRHQX1 \funct_out_reg[1]  ( .D(funct_in[1]), .CK(clk), .RN(rst), .Q(
        funct_out[1]) );
  DFFRHQX1 \funct_out_reg[2]  ( .D(funct_in[2]), .CK(clk), .RN(rst), .Q(
        funct_out[2]) );
  DFFRHQX1 \read_data1_out_reg[21]  ( .D(read_data1_in[21]), .CK(clk), .RN(rst), .Q(read_data1_out[21]) );
  DFFRHQX1 \read_data1_out_reg[20]  ( .D(read_data1_in[20]), .CK(clk), .RN(rst), .Q(read_data1_out[20]) );
  DFFRHQX1 \read_data1_out_reg[19]  ( .D(read_data1_in[19]), .CK(clk), .RN(rst), .Q(read_data1_out[19]) );
  DFFRHQX1 \read_data1_out_reg[18]  ( .D(read_data1_in[18]), .CK(clk), .RN(rst), .Q(read_data1_out[18]) );
  DFFRHQX1 \read_data1_out_reg[17]  ( .D(read_data1_in[17]), .CK(clk), .RN(rst), .Q(read_data1_out[17]) );
  DFFRHQX1 \read_data1_out_reg[16]  ( .D(read_data1_in[16]), .CK(clk), .RN(rst), .Q(read_data1_out[16]) );
  DFFRHQX1 \read_data1_out_reg[15]  ( .D(read_data1_in[15]), .CK(clk), .RN(rst), .Q(read_data1_out[15]) );
  DFFRHQX1 \read_data1_out_reg[14]  ( .D(read_data1_in[14]), .CK(clk), .RN(rst), .Q(read_data1_out[14]) );
  DFFRHQX1 \read_data1_out_reg[13]  ( .D(read_data1_in[13]), .CK(clk), .RN(rst), .Q(read_data1_out[13]) );
  DFFRHQX1 \read_data1_out_reg[12]  ( .D(read_data1_in[12]), .CK(clk), .RN(rst), .Q(read_data1_out[12]) );
  DFFRHQX1 \read_data1_out_reg[11]  ( .D(read_data1_in[11]), .CK(clk), .RN(rst), .Q(read_data1_out[11]) );
  DFFRHQX1 \read_data2_out_reg[31]  ( .D(read_data2_in[31]), .CK(clk), .RN(rst), .Q(read_data2_out[31]) );
  DFFRHQX1 \read_data2_out_reg[30]  ( .D(read_data2_in[30]), .CK(clk), .RN(rst), .Q(read_data2_out[30]) );
  DFFRHQX1 \read_data2_out_reg[29]  ( .D(read_data2_in[29]), .CK(clk), .RN(rst), .Q(read_data2_out[29]) );
  DFFRHQX1 \read_data2_out_reg[28]  ( .D(read_data2_in[28]), .CK(clk), .RN(rst), .Q(read_data2_out[28]) );
  DFFRHQX1 \read_data2_out_reg[27]  ( .D(read_data2_in[27]), .CK(clk), .RN(rst), .Q(read_data2_out[27]) );
  DFFRHQX1 \read_data2_out_reg[26]  ( .D(read_data2_in[26]), .CK(clk), .RN(rst), .Q(read_data2_out[26]) );
  DFFRHQX1 \read_data2_out_reg[25]  ( .D(read_data2_in[25]), .CK(clk), .RN(rst), .Q(read_data2_out[25]) );
  DFFRHQX1 \read_data2_out_reg[24]  ( .D(read_data2_in[24]), .CK(clk), .RN(rst), .Q(read_data2_out[24]) );
  DFFRHQX1 \read_data2_out_reg[23]  ( .D(read_data2_in[23]), .CK(clk), .RN(rst), .Q(read_data2_out[23]) );
  DFFRHQX1 \read_data2_out_reg[22]  ( .D(read_data2_in[22]), .CK(clk), .RN(rst), .Q(read_data2_out[22]) );
  DFFRHQX1 \read_data2_out_reg[21]  ( .D(read_data2_in[21]), .CK(clk), .RN(rst), .Q(read_data2_out[21]) );
  DFFRHQX1 \read_data2_out_reg[20]  ( .D(read_data2_in[20]), .CK(clk), .RN(rst), .Q(read_data2_out[20]) );
  DFFRHQX1 \read_data2_out_reg[19]  ( .D(read_data2_in[19]), .CK(clk), .RN(rst), .Q(read_data2_out[19]) );
  DFFRHQX1 \read_data2_out_reg[18]  ( .D(read_data2_in[18]), .CK(clk), .RN(rst), .Q(read_data2_out[18]) );
  DFFRHQX1 \read_data2_out_reg[17]  ( .D(read_data2_in[17]), .CK(clk), .RN(rst), .Q(read_data2_out[17]) );
  DFFRHQX1 \read_data2_out_reg[16]  ( .D(read_data2_in[16]), .CK(clk), .RN(rst), .Q(read_data2_out[16]) );
  DFFRHQX1 \read_data2_out_reg[15]  ( .D(read_data2_in[15]), .CK(clk), .RN(rst), .Q(read_data2_out[15]) );
  DFFRHQX1 \read_data2_out_reg[14]  ( .D(read_data2_in[14]), .CK(clk), .RN(rst), .Q(read_data2_out[14]) );
  DFFRHQX1 \read_data2_out_reg[13]  ( .D(read_data2_in[13]), .CK(clk), .RN(rst), .Q(read_data2_out[13]) );
  DFFRHQX1 \ext_out_reg[31]  ( .D(ext_in[31]), .CK(clk), .RN(rst), .Q(
        ext_out[31]) );
  DFFRHQX1 \ext_out_reg[30]  ( .D(ext_in[30]), .CK(clk), .RN(rst), .Q(
        ext_out[30]) );
  DFFRHQX1 \ext_out_reg[29]  ( .D(ext_in[29]), .CK(clk), .RN(rst), .Q(
        ext_out[29]) );
  DFFRHQX1 \ext_out_reg[28]  ( .D(ext_in[28]), .CK(clk), .RN(rst), .Q(
        ext_out[28]) );
  DFFRHQX1 \ext_out_reg[27]  ( .D(ext_in[27]), .CK(clk), .RN(rst), .Q(
        ext_out[27]) );
  DFFRHQX1 \ext_out_reg[26]  ( .D(ext_in[26]), .CK(clk), .RN(rst), .Q(
        ext_out[26]) );
  DFFRHQX1 \ext_out_reg[25]  ( .D(ext_in[25]), .CK(clk), .RN(rst), .Q(
        ext_out[25]) );
  DFFRHQX1 \ext_out_reg[24]  ( .D(ext_in[24]), .CK(clk), .RN(rst), .Q(
        ext_out[24]) );
  DFFRHQX1 \ext_out_reg[23]  ( .D(ext_in[23]), .CK(clk), .RN(rst), .Q(
        ext_out[23]) );
  DFFRHQX1 \ext_out_reg[22]  ( .D(ext_in[22]), .CK(clk), .RN(rst), .Q(
        ext_out[22]) );
  DFFRHQX1 \ext_out_reg[21]  ( .D(ext_in[21]), .CK(clk), .RN(rst), .Q(
        ext_out[21]) );
  DFFRHQX1 \ext_out_reg[20]  ( .D(ext_in[20]), .CK(clk), .RN(rst), .Q(
        ext_out[20]) );
  DFFRHQX1 \ext_out_reg[19]  ( .D(ext_in[19]), .CK(clk), .RN(rst), .Q(
        ext_out[19]) );
  DFFRHQX1 \ext_out_reg[18]  ( .D(ext_in[18]), .CK(clk), .RN(rst), .Q(
        ext_out[18]) );
  DFFRHQX1 \ext_out_reg[17]  ( .D(ext_in[17]), .CK(clk), .RN(rst), .Q(
        ext_out[17]) );
  DFFRHQX1 \ext_out_reg[16]  ( .D(ext_in[16]), .CK(clk), .RN(rst), .Q(
        ext_out[16]) );
  DFFRHQX1 \ext_out_reg[15]  ( .D(ext_in[15]), .CK(clk), .RN(rst), .Q(
        ext_out[15]) );
  DFFRHQX1 \ext_out_reg[14]  ( .D(ext_in[14]), .CK(clk), .RN(rst), .Q(
        ext_out[14]) );
  DFFRHQX1 \ext_out_reg[13]  ( .D(ext_in[13]), .CK(clk), .RN(rst), .Q(
        ext_out[13]) );
  DFFRHQX1 \read_data1_out_reg[10]  ( .D(read_data1_in[10]), .CK(clk), .RN(rst), .Q(read_data1_out[10]) );
  DFFRHQX1 \read_data1_out_reg[9]  ( .D(read_data1_in[9]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[9]) );
  DFFRHQX1 \read_data1_out_reg[8]  ( .D(read_data1_in[8]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[8]) );
  DFFRHQX1 \read_data1_out_reg[7]  ( .D(read_data1_in[7]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[7]) );
  DFFRHQX1 \read_data1_out_reg[6]  ( .D(read_data1_in[6]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[6]) );
  DFFRHQX1 \read_data1_out_reg[5]  ( .D(read_data1_in[5]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[5]) );
  DFFRHQX1 \read_data1_out_reg[4]  ( .D(read_data1_in[4]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[4]) );
  DFFRHQX1 \read_data1_out_reg[3]  ( .D(read_data1_in[3]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[3]) );
  DFFRHQX1 \read_data1_out_reg[2]  ( .D(read_data1_in[2]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[2]) );
  DFFRHQX1 \read_data1_out_reg[1]  ( .D(read_data1_in[1]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[1]) );
  DFFRHQX1 \read_data1_out_reg[0]  ( .D(read_data1_in[0]), .CK(clk), .RN(rst), 
        .Q(read_data1_out[0]) );
  DFFRHQX1 \read_data2_out_reg[12]  ( .D(read_data2_in[12]), .CK(clk), .RN(rst), .Q(read_data2_out[12]) );
  DFFRHQX1 \read_data2_out_reg[11]  ( .D(read_data2_in[11]), .CK(clk), .RN(rst), .Q(read_data2_out[11]) );
  DFFRHQX1 \read_data2_out_reg[10]  ( .D(read_data2_in[10]), .CK(clk), .RN(rst), .Q(read_data2_out[10]) );
  DFFRHQX1 \read_data2_out_reg[9]  ( .D(read_data2_in[9]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[9]) );
  DFFRHQX1 \read_data2_out_reg[8]  ( .D(read_data2_in[8]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[8]) );
  DFFRHQX1 \read_data2_out_reg[7]  ( .D(read_data2_in[7]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[7]) );
  DFFRHQX1 \read_data2_out_reg[6]  ( .D(read_data2_in[6]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[6]) );
  DFFRHQX1 \read_data2_out_reg[5]  ( .D(read_data2_in[5]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[5]) );
  DFFRHQX1 \read_data2_out_reg[4]  ( .D(read_data2_in[4]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[4]) );
  DFFRHQX1 \read_data2_out_reg[3]  ( .D(read_data2_in[3]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[3]) );
  DFFRHQX1 \read_data2_out_reg[2]  ( .D(read_data2_in[2]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[2]) );
  DFFRHQX1 \ext_out_reg[12]  ( .D(ext_in[12]), .CK(clk), .RN(rst), .Q(
        ext_out[12]) );
  DFFRHQX1 \ext_out_reg[11]  ( .D(ext_in[11]), .CK(clk), .RN(rst), .Q(
        ext_out[11]) );
  DFFRHQX1 \ext_out_reg[10]  ( .D(ext_in[10]), .CK(clk), .RN(rst), .Q(
        ext_out[10]) );
  DFFRHQX1 \ext_out_reg[8]  ( .D(ext_in[8]), .CK(clk), .RN(rst), .Q(ext_out[8]) );
  DFFRHQX1 \ext_out_reg[7]  ( .D(ext_in[7]), .CK(clk), .RN(rst), .Q(ext_out[7]) );
  DFFRHQX1 \ext_out_reg[6]  ( .D(ext_in[6]), .CK(clk), .RN(rst), .Q(ext_out[6]) );
  DFFRHQX1 \ext_out_reg[5]  ( .D(ext_in[5]), .CK(clk), .RN(rst), .Q(ext_out[5]) );
  DFFRHQX1 \ext_out_reg[4]  ( .D(ext_in[4]), .CK(clk), .RN(rst), .Q(ext_out[4]) );
  DFFRHQX1 \ext_out_reg[3]  ( .D(ext_in[3]), .CK(clk), .RN(rst), .Q(ext_out[3]) );
  DFFRHQX1 \ext_out_reg[2]  ( .D(ext_in[2]), .CK(clk), .RN(rst), .Q(ext_out[2]) );
  DFFRHQX1 \ext_out_reg[9]  ( .D(ext_in[9]), .CK(clk), .RN(rst), .Q(ext_out[9]) );
  DFFRHQX1 \inst_out_reg[8]  ( .D(inst_in[8]), .CK(clk), .RN(rst), .Q(
        inst_out[8]) );
  DFFRHQX1 \inst_out_reg[9]  ( .D(inst_in[9]), .CK(clk), .RN(rst), .Q(
        inst_out[9]) );
  DFFRHQX1 \addr1_out_reg[3]  ( .D(addr1_in[3]), .CK(clk), .RN(rst), .Q(
        addr1_out[3]) );
  DFFRHQX1 \addr2_out_reg[3]  ( .D(addr2_in[3]), .CK(clk), .RN(rst), .Q(
        addr2_out[3]) );
  DFFRHQX1 \addr1_out_reg[4]  ( .D(addr1_in[4]), .CK(clk), .RN(rst), .Q(
        addr1_out[4]) );
  DFFRHQX1 \addr1_out_reg[2]  ( .D(addr1_in[2]), .CK(clk), .RN(rst), .Q(
        addr1_out[2]) );
  DFFRHQX1 \addr1_out_reg[0]  ( .D(addr1_in[0]), .CK(clk), .RN(rst), .Q(
        addr1_out[0]) );
  DFFRHQX1 \addr2_out_reg[4]  ( .D(addr2_in[4]), .CK(clk), .RN(rst), .Q(
        addr2_out[4]) );
  DFFRHQX1 \addr2_out_reg[2]  ( .D(addr2_in[2]), .CK(clk), .RN(rst), .Q(
        addr2_out[2]) );
  DFFRHQX1 \addr2_out_reg[0]  ( .D(addr2_in[0]), .CK(clk), .RN(rst), .Q(
        addr2_out[0]) );
  DFFRHQX1 \addr1_out_reg[1]  ( .D(addr1_in[1]), .CK(clk), .RN(rst), .Q(
        addr1_out[1]) );
  DFFRHQX1 \addr2_out_reg[1]  ( .D(addr2_in[1]), .CK(clk), .RN(rst), .Q(
        addr2_out[1]) );
  DFFRHQX1 \read_data2_out_reg[1]  ( .D(read_data2_in[1]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[1]) );
  DFFRHQX1 \read_data2_out_reg[0]  ( .D(read_data2_in[0]), .CK(clk), .RN(rst), 
        .Q(read_data2_out[0]) );
  DFFRHQX1 ls_w_mode_out_reg ( .D(ls_w_mode_in), .CK(clk), .RN(rst), .Q(
        ls_w_mode_out) );
  DFFRHQX1 \ext_out_reg[1]  ( .D(ext_in[1]), .CK(clk), .RN(rst), .Q(ext_out[1]) );
  DFFRHQX1 \ext_out_reg[0]  ( .D(ext_in[0]), .CK(clk), .RN(rst), .Q(ext_out[0]) );
  DFFRHQX1 sel_in2_out_reg ( .D(sel_in2_in), .CK(clk), .RN(rst), .Q(
        sel_in2_out) );
  DFFRHQX1 \inst_out_reg[24]  ( .D(inst_in[24]), .CK(clk), .RN(rst), .Q(
        inst_out[24]) );
  DFFRHQX1 \inst_out_reg[23]  ( .D(inst_in[23]), .CK(clk), .RN(rst), .Q(
        inst_out[23]) );
  DFFRHQX1 \inst_out_reg[22]  ( .D(inst_in[22]), .CK(clk), .RN(rst), .Q(
        inst_out[22]) );
  DFFRHQX1 \inst_out_reg[21]  ( .D(inst_in[21]), .CK(clk), .RN(rst), .Q(
        inst_out[21]) );
  DFFRHQX1 \inst_out_reg[20]  ( .D(inst_in[20]), .CK(clk), .RN(rst), .Q(
        inst_out[20]) );
  DFFRHQX1 \inst_out_reg[19]  ( .D(inst_in[19]), .CK(clk), .RN(rst), .Q(
        inst_out[19]) );
  DFFRHQX1 \inst_out_reg[18]  ( .D(inst_in[18]), .CK(clk), .RN(rst), .Q(
        inst_out[18]) );
  DFFRHQX1 \inst_out_reg[17]  ( .D(inst_in[17]), .CK(clk), .RN(rst), .Q(
        inst_out[17]) );
  DFFRHQX1 \inst_out_reg[16]  ( .D(inst_in[16]), .CK(clk), .RN(rst), .Q(
        inst_out[16]) );
  DFFRHQX1 \inst_out_reg[15]  ( .D(inst_in[15]), .CK(clk), .RN(rst), .Q(
        inst_out[15]) );
  DFFRHQX1 \inst_out_reg[14]  ( .D(inst_in[14]), .CK(clk), .RN(rst), .Q(
        inst_out[14]) );
  DFFRHQX1 \inst_out_reg[13]  ( .D(inst_in[13]), .CK(clk), .RN(rst), .Q(
        inst_out[13]) );
  DFFRHQX1 \inst_out_reg[12]  ( .D(inst_in[12]), .CK(clk), .RN(rst), .Q(
        inst_out[12]) );
  DFFRHQX1 \inst_out_reg[11]  ( .D(inst_in[11]), .CK(clk), .RN(rst), .Q(
        inst_out[11]) );
  DFFRHQX1 \inst_out_reg[10]  ( .D(inst_in[10]), .CK(clk), .RN(rst), .Q(
        inst_out[10]) );
  DFFRHQX1 \read_data3_out_reg[31]  ( .D(read_data3_in[31]), .CK(clk), .RN(rst), .Q(read_data3_out[31]) );
  DFFRHQX1 \read_data3_out_reg[30]  ( .D(read_data3_in[30]), .CK(clk), .RN(rst), .Q(read_data3_out[30]) );
  DFFRHQX1 \read_data3_out_reg[29]  ( .D(read_data3_in[29]), .CK(clk), .RN(rst), .Q(read_data3_out[29]) );
  DFFRHQX1 \read_data3_out_reg[28]  ( .D(read_data3_in[28]), .CK(clk), .RN(rst), .Q(read_data3_out[28]) );
  DFFRHQX1 \read_data3_out_reg[27]  ( .D(read_data3_in[27]), .CK(clk), .RN(rst), .Q(read_data3_out[27]) );
  DFFRHQX1 \read_data3_out_reg[26]  ( .D(read_data3_in[26]), .CK(clk), .RN(rst), .Q(read_data3_out[26]) );
  DFFRHQX1 \read_data3_out_reg[25]  ( .D(read_data3_in[25]), .CK(clk), .RN(rst), .Q(read_data3_out[25]) );
  DFFRHQX1 \read_data3_out_reg[24]  ( .D(read_data3_in[24]), .CK(clk), .RN(rst), .Q(read_data3_out[24]) );
  DFFRHQX1 \read_data3_out_reg[23]  ( .D(read_data3_in[23]), .CK(clk), .RN(rst), .Q(read_data3_out[23]) );
  DFFRHQX1 \read_data3_out_reg[22]  ( .D(read_data3_in[22]), .CK(clk), .RN(rst), .Q(read_data3_out[22]) );
  DFFRHQX1 \read_data3_out_reg[21]  ( .D(read_data3_in[21]), .CK(clk), .RN(rst), .Q(read_data3_out[21]) );
  DFFRHQX1 \read_data3_out_reg[20]  ( .D(read_data3_in[20]), .CK(clk), .RN(rst), .Q(read_data3_out[20]) );
  DFFRHQX1 \read_data3_out_reg[19]  ( .D(read_data3_in[19]), .CK(clk), .RN(rst), .Q(read_data3_out[19]) );
  DFFRHQX1 \read_data3_out_reg[18]  ( .D(read_data3_in[18]), .CK(clk), .RN(rst), .Q(read_data3_out[18]) );
  DFFRHQX1 \read_data3_out_reg[17]  ( .D(read_data3_in[17]), .CK(clk), .RN(rst), .Q(read_data3_out[17]) );
  DFFRHQX1 \read_data3_out_reg[16]  ( .D(read_data3_in[16]), .CK(clk), .RN(rst), .Q(read_data3_out[16]) );
  DFFRHQX1 \read_data3_out_reg[15]  ( .D(read_data3_in[15]), .CK(clk), .RN(rst), .Q(read_data3_out[15]) );
  DFFRHQX1 \read_data3_out_reg[14]  ( .D(read_data3_in[14]), .CK(clk), .RN(rst), .Q(read_data3_out[14]) );
  DFFRHQX1 \read_data3_out_reg[13]  ( .D(read_data3_in[13]), .CK(clk), .RN(rst), .Q(read_data3_out[13]) );
  DFFRHQX1 \read_data3_out_reg[12]  ( .D(read_data3_in[12]), .CK(clk), .RN(rst), .Q(read_data3_out[12]) );
  DFFRHQX1 \read_data3_out_reg[11]  ( .D(read_data3_in[11]), .CK(clk), .RN(rst), .Q(read_data3_out[11]) );
  DFFRHQX1 \read_data3_out_reg[10]  ( .D(read_data3_in[10]), .CK(clk), .RN(rst), .Q(read_data3_out[10]) );
  DFFRHQX1 \read_data3_out_reg[9]  ( .D(read_data3_in[9]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[9]) );
  DFFRHQX1 \read_data3_out_reg[8]  ( .D(read_data3_in[8]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[8]) );
  DFFRHQX1 \read_data3_out_reg[7]  ( .D(read_data3_in[7]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[7]) );
  DFFRHQX1 \read_data3_out_reg[6]  ( .D(read_data3_in[6]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[6]) );
  DFFRHQX1 \read_data3_out_reg[5]  ( .D(read_data3_in[5]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[5]) );
  DFFRHQX1 \read_data3_out_reg[4]  ( .D(read_data3_in[4]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[4]) );
  DFFRHQX1 \read_data3_out_reg[3]  ( .D(read_data3_in[3]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[3]) );
  DFFRHQX1 \read_data3_out_reg[2]  ( .D(read_data3_in[2]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[2]) );
  DFFRHQX1 \read_data3_out_reg[1]  ( .D(read_data3_in[1]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[1]) );
  DFFRHQX1 \read_data3_out_reg[0]  ( .D(read_data3_in[0]), .CK(clk), .RN(rst), 
        .Q(read_data3_out[0]) );
  DFFRHQX1 data_rw_out_reg ( .D(data_rw_in), .CK(clk), .RN(rst), .Q(
        data_rw_out) );
  DFFRHQX1 sel_wb_out_reg ( .D(sel_wb_in), .CK(clk), .RN(rst), .Q(sel_wb_out)
         );
  DFFRHQX1 reg_rw_out_reg ( .D(reg_rw_in), .CK(clk), .RN(rst), .Q(reg_rw_out)
         );
  DFFRHQX1 \inst_out_reg[31]  ( .D(inst_in[31]), .CK(clk), .RN(rst), .Q(
        inst_out[31]) );
  DFFRHQX1 \inst_out_reg[30]  ( .D(inst_in[30]), .CK(clk), .RN(rst), .Q(
        inst_out[30]) );
  DFFRHQX1 \inst_out_reg[29]  ( .D(inst_in[29]), .CK(clk), .RN(rst), .Q(
        inst_out[29]) );
  DFFRHQX1 \inst_out_reg[28]  ( .D(inst_in[28]), .CK(clk), .RN(rst), .Q(
        inst_out[28]) );
  DFFRHQX1 \inst_out_reg[27]  ( .D(inst_in[27]), .CK(clk), .RN(rst), .Q(
        inst_out[27]) );
  DFFRHQX1 \inst_out_reg[26]  ( .D(inst_in[26]), .CK(clk), .RN(rst), .Q(
        inst_out[26]) );
  DFFRHQX1 \inst_out_reg[25]  ( .D(inst_in[25]), .CK(clk), .RN(rst), .Q(
        inst_out[25]) );
  DFFRHQX1 \inst_out_reg[7]  ( .D(inst_in[7]), .CK(clk), .RN(rst), .Q(
        inst_out[7]) );
  DFFRHQX1 \inst_out_reg[6]  ( .D(inst_in[6]), .CK(clk), .RN(rst), .Q(
        inst_out[6]) );
  DFFRHQX1 \inst_out_reg[5]  ( .D(inst_in[5]), .CK(clk), .RN(rst), .Q(
        inst_out[5]) );
  DFFRHQX1 \inst_out_reg[4]  ( .D(inst_in[4]), .CK(clk), .RN(rst), .Q(
        inst_out[4]) );
  DFFRHQX1 \inst_out_reg[3]  ( .D(inst_in[3]), .CK(clk), .RN(rst), .Q(
        inst_out[3]) );
  DFFRHQX1 \inst_out_reg[2]  ( .D(inst_in[2]), .CK(clk), .RN(rst), .Q(
        inst_out[2]) );
  DFFRHQX1 \inst_out_reg[1]  ( .D(inst_in[1]), .CK(clk), .RN(rst), .Q(
        inst_out[1]) );
  DFFRHQX1 \inst_out_reg[0]  ( .D(inst_in[0]), .CK(clk), .RN(rst), .Q(
        inst_out[0]) );
endmodule


module CONTROLLER ( reg_ena, funct, ls_w_mode, sign_ena, sel_in2, ena_data, 
        data_rw, sel_wb, reg_rw, sel, opcode, subopcode, read_data1, 
        read_data2, clk, rst, sel_alu, branch_ena, Jump_ena );
  output [3:0] funct;
  output [2:0] sel;
  input [5:0] opcode;
  input [4:0] subopcode;
  input [31:0] read_data1;
  input [31:0] read_data2;
  input clk, rst;
  output reg_ena, ls_w_mode, sign_ena, sel_in2, ena_data, data_rw, sel_wb,
         reg_rw, sel_alu, branch_ena, Jump_ena;
  wire   Jump_ena, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49;
  assign reg_ena = 1'b1;
  assign sel[2] = Jump_ena;

  INVX1 U3 ( .A(n15), .Y(Jump_ena) );
  INVX1 U4 ( .A(n14), .Y(sel[0]) );
  OR2X2 U5 ( .A(ena_data), .B(sel_wb), .Y(reg_rw) );
  NAND3X1 U6 ( .A(n24), .B(n25), .C(n26), .Y(sel[1]) );
  NOR2X1 U7 ( .A(branch_ena), .B(sel_alu), .Y(n14) );
  NAND2X1 U8 ( .A(n22), .B(n23), .Y(n15) );
  AND4X2 U9 ( .A(n32), .B(n33), .C(n28), .D(n13), .Y(n26) );
  INVX1 U10 ( .A(n25), .Y(sel_alu) );
  NAND3X1 U11 ( .A(n13), .B(n14), .C(n15), .Y(sign_ena) );
  NAND3X1 U12 ( .A(n45), .B(n29), .C(n23), .Y(n21) );
  INVX1 U13 ( .A(n18), .Y(n34) );
  OAI21XL U14 ( .A0(n49), .A1(n30), .B0(n32), .Y(data_rw) );
  OAI33X1 U15 ( .A0(n16), .A1(n17), .A2(n18), .B0(n19), .B1(n20), .B2(
        ls_w_mode), .Y(sel_in2) );
  INVX1 U16 ( .A(n21), .Y(n20) );
  NAND2X1 U17 ( .A(n15), .B(n14), .Y(n19) );
  NAND4X1 U18 ( .A(n26), .B(n43), .C(n30), .D(n35), .Y(funct[0]) );
  NAND3X1 U19 ( .A(n41), .B(n16), .C(n34), .Y(n43) );
  OAI221XL U20 ( .A0(n18), .A1(n41), .B0(n21), .B1(n42), .C0(n35), .Y(funct[1]) );
  OAI21XL U21 ( .A0(n42), .A1(n30), .B0(n33), .Y(ena_data) );
  NAND4X1 U22 ( .A(n13), .B(n25), .C(n21), .D(n27), .Y(sel_wb) );
  AND2X2 U23 ( .A(n24), .B(n28), .Y(n27) );
  INVX1 U24 ( .A(n49), .Y(n42) );
  INVX1 U25 ( .A(n30), .Y(ls_w_mode) );
  NOR3X1 U26 ( .A(opcode[2]), .B(opcode[4]), .C(n45), .Y(n47) );
  AND3X2 U27 ( .A(opcode[1]), .B(n23), .C(opcode[2]), .Y(branch_ena) );
  NOR3BX1 U28 ( .AN(opcode[5]), .B(opcode[0]), .C(opcode[4]), .Y(n40) );
  NAND3X1 U29 ( .A(n23), .B(n29), .C(opcode[1]), .Y(n25) );
  NOR2BX1 U30 ( .AN(n40), .B(opcode[3]), .Y(n23) );
  NOR2X1 U31 ( .A(n29), .B(opcode[1]), .Y(n22) );
  NAND4X1 U32 ( .A(opcode[3]), .B(n40), .C(n45), .D(n29), .Y(n13) );
  NOR2X1 U33 ( .A(opcode[5]), .B(opcode[0]), .Y(n48) );
  NAND3BX1 U34 ( .AN(opcode[3]), .B(n47), .C(n48), .Y(n33) );
  NAND3X1 U35 ( .A(n47), .B(opcode[3]), .C(n48), .Y(n32) );
  NAND4X1 U36 ( .A(opcode[0]), .B(n47), .C(opcode[3]), .D(opcode[5]), .Y(n28)
         );
  INVX1 U37 ( .A(opcode[2]), .Y(n29) );
  INVX1 U38 ( .A(opcode[1]), .Y(n45) );
  NAND3X1 U39 ( .A(opcode[3]), .B(n40), .C(n22), .Y(n24) );
  NOR2X1 U40 ( .A(n21), .B(subopcode[4]), .Y(n37) );
  NAND2BX1 U41 ( .AN(subopcode[2]), .B(n37), .Y(n18) );
  NAND4X1 U42 ( .A(n24), .B(n35), .C(n28), .D(n36), .Y(funct[2]) );
  AOI33X1 U43 ( .A0(subopcode[2]), .A1(n37), .A2(n38), .B0(n34), .B1(n39), 
        .B2(subopcode[0]), .Y(n36) );
  NOR3X1 U44 ( .A(subopcode[0]), .B(subopcode[3]), .C(subopcode[1]), .Y(n38)
         );
  NAND4X1 U45 ( .A(n31), .B(n32), .C(n33), .D(n30), .Y(funct[3]) );
  NAND4X1 U46 ( .A(subopcode[0]), .B(subopcode[3]), .C(n34), .D(subopcode[1]), 
        .Y(n31) );
  NOR4BX1 U47 ( .AN(n17), .B(subopcode[2]), .C(subopcode[3]), .D(subopcode[4]), 
        .Y(n49) );
  NAND4X1 U48 ( .A(opcode[4]), .B(n48), .C(n22), .D(opcode[3]), .Y(n30) );
  NAND3X1 U49 ( .A(subopcode[3]), .B(n37), .C(n44), .Y(n35) );
  NOR3X1 U50 ( .A(subopcode[0]), .B(subopcode[2]), .C(subopcode[1]), .Y(n44)
         );
  NAND2X1 U51 ( .A(subopcode[0]), .B(n46), .Y(n41) );
  NOR2X1 U52 ( .A(n46), .B(subopcode[0]), .Y(n17) );
  INVX1 U53 ( .A(subopcode[1]), .Y(n46) );
  INVX1 U54 ( .A(subopcode[3]), .Y(n16) );
  XNOR2X1 U55 ( .A(n16), .B(subopcode[1]), .Y(n39) );
endmodule


module REGISTER_FILE ( clk, rst, reg_rw, reg_ena, addr1, addr2, addr_dst, 
        write_data, write_addr, read_data1, read_data2, read_data3 );
  input [4:0] addr1;
  input [4:0] addr2;
  input [4:0] addr_dst;
  input [31:0] write_data;
  input [4:0] write_addr;
  output [31:0] read_data1;
  output [31:0] read_data2;
  output [31:0] read_data3;
  input clk, rst, reg_rw, reg_ena;
  wire   N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, \regs[31][31] , \regs[31][30] , \regs[31][29] , \regs[31][28] ,
         \regs[31][27] , \regs[31][26] , \regs[31][25] , \regs[31][24] ,
         \regs[31][23] , \regs[31][22] , \regs[31][21] , \regs[31][20] ,
         \regs[31][19] , \regs[31][18] , \regs[31][17] , \regs[31][16] ,
         \regs[31][15] , \regs[31][14] , \regs[31][13] , \regs[31][12] ,
         \regs[31][11] , \regs[31][10] , \regs[31][9] , \regs[31][8] ,
         \regs[31][7] , \regs[31][6] , \regs[31][5] , \regs[31][4] ,
         \regs[31][3] , \regs[31][2] , \regs[31][1] , \regs[31][0] ,
         \regs[30][31] , \regs[30][30] , \regs[30][29] , \regs[30][28] ,
         \regs[30][27] , \regs[30][26] , \regs[30][25] , \regs[30][24] ,
         \regs[30][23] , \regs[30][22] , \regs[30][21] , \regs[30][20] ,
         \regs[30][19] , \regs[30][18] , \regs[30][17] , \regs[30][16] ,
         \regs[30][15] , \regs[30][14] , \regs[30][13] , \regs[30][12] ,
         \regs[30][11] , \regs[30][10] , \regs[30][9] , \regs[30][8] ,
         \regs[30][7] , \regs[30][6] , \regs[30][5] , \regs[30][4] ,
         \regs[30][3] , \regs[30][2] , \regs[30][1] , \regs[30][0] ,
         \regs[29][31] , \regs[29][30] , \regs[29][29] , \regs[29][28] ,
         \regs[29][27] , \regs[29][26] , \regs[29][25] , \regs[29][24] ,
         \regs[29][23] , \regs[29][22] , \regs[29][21] , \regs[29][20] ,
         \regs[29][19] , \regs[29][18] , \regs[29][17] , \regs[29][16] ,
         \regs[29][15] , \regs[29][14] , \regs[29][13] , \regs[29][12] ,
         \regs[29][11] , \regs[29][10] , \regs[29][9] , \regs[29][8] ,
         \regs[29][7] , \regs[29][6] , \regs[29][5] , \regs[29][4] ,
         \regs[29][3] , \regs[29][2] , \regs[29][1] , \regs[29][0] ,
         \regs[28][31] , \regs[28][30] , \regs[28][29] , \regs[28][28] ,
         \regs[28][27] , \regs[28][26] , \regs[28][25] , \regs[28][24] ,
         \regs[28][23] , \regs[28][22] , \regs[28][21] , \regs[28][20] ,
         \regs[28][19] , \regs[28][18] , \regs[28][17] , \regs[28][16] ,
         \regs[28][15] , \regs[28][14] , \regs[28][13] , \regs[28][12] ,
         \regs[28][11] , \regs[28][10] , \regs[28][9] , \regs[28][8] ,
         \regs[28][7] , \regs[28][6] , \regs[28][5] , \regs[28][4] ,
         \regs[28][3] , \regs[28][2] , \regs[28][1] , \regs[28][0] ,
         \regs[27][31] , \regs[27][30] , \regs[27][29] , \regs[27][28] ,
         \regs[27][27] , \regs[27][26] , \regs[27][25] , \regs[27][24] ,
         \regs[27][23] , \regs[27][22] , \regs[27][21] , \regs[27][20] ,
         \regs[27][19] , \regs[27][18] , \regs[27][17] , \regs[27][16] ,
         \regs[27][15] , \regs[27][14] , \regs[27][13] , \regs[27][12] ,
         \regs[27][11] , \regs[27][10] , \regs[27][9] , \regs[27][8] ,
         \regs[27][7] , \regs[27][6] , \regs[27][5] , \regs[27][4] ,
         \regs[27][3] , \regs[27][2] , \regs[27][1] , \regs[27][0] ,
         \regs[26][31] , \regs[26][30] , \regs[26][29] , \regs[26][28] ,
         \regs[26][27] , \regs[26][26] , \regs[26][25] , \regs[26][24] ,
         \regs[26][23] , \regs[26][22] , \regs[26][21] , \regs[26][20] ,
         \regs[26][19] , \regs[26][18] , \regs[26][17] , \regs[26][16] ,
         \regs[26][15] , \regs[26][14] , \regs[26][13] , \regs[26][12] ,
         \regs[26][11] , \regs[26][10] , \regs[26][9] , \regs[26][8] ,
         \regs[26][7] , \regs[26][6] , \regs[26][5] , \regs[26][4] ,
         \regs[26][3] , \regs[26][2] , \regs[26][1] , \regs[26][0] ,
         \regs[25][31] , \regs[25][30] , \regs[25][29] , \regs[25][28] ,
         \regs[25][27] , \regs[25][26] , \regs[25][25] , \regs[25][24] ,
         \regs[25][23] , \regs[25][22] , \regs[25][21] , \regs[25][20] ,
         \regs[25][19] , \regs[25][18] , \regs[25][17] , \regs[25][16] ,
         \regs[25][15] , \regs[25][14] , \regs[25][13] , \regs[25][12] ,
         \regs[25][11] , \regs[25][10] , \regs[25][9] , \regs[25][8] ,
         \regs[25][7] , \regs[25][6] , \regs[25][5] , \regs[25][4] ,
         \regs[25][3] , \regs[25][2] , \regs[25][1] , \regs[25][0] ,
         \regs[24][31] , \regs[24][30] , \regs[24][29] , \regs[24][28] ,
         \regs[24][27] , \regs[24][26] , \regs[24][25] , \regs[24][24] ,
         \regs[24][23] , \regs[24][22] , \regs[24][21] , \regs[24][20] ,
         \regs[24][19] , \regs[24][18] , \regs[24][17] , \regs[24][16] ,
         \regs[24][15] , \regs[24][14] , \regs[24][13] , \regs[24][12] ,
         \regs[24][11] , \regs[24][10] , \regs[24][9] , \regs[24][8] ,
         \regs[24][7] , \regs[24][6] , \regs[24][5] , \regs[24][4] ,
         \regs[24][3] , \regs[24][2] , \regs[24][1] , \regs[24][0] ,
         \regs[23][31] , \regs[23][30] , \regs[23][29] , \regs[23][28] ,
         \regs[23][27] , \regs[23][26] , \regs[23][25] , \regs[23][24] ,
         \regs[23][23] , \regs[23][22] , \regs[23][21] , \regs[23][20] ,
         \regs[23][19] , \regs[23][18] , \regs[23][17] , \regs[23][16] ,
         \regs[23][15] , \regs[23][14] , \regs[23][13] , \regs[23][12] ,
         \regs[23][11] , \regs[23][10] , \regs[23][9] , \regs[23][8] ,
         \regs[23][7] , \regs[23][6] , \regs[23][5] , \regs[23][4] ,
         \regs[23][3] , \regs[23][2] , \regs[23][1] , \regs[23][0] ,
         \regs[22][31] , \regs[22][30] , \regs[22][29] , \regs[22][28] ,
         \regs[22][27] , \regs[22][26] , \regs[22][25] , \regs[22][24] ,
         \regs[22][23] , \regs[22][22] , \regs[22][21] , \regs[22][20] ,
         \regs[22][19] , \regs[22][18] , \regs[22][17] , \regs[22][16] ,
         \regs[22][15] , \regs[22][14] , \regs[22][13] , \regs[22][12] ,
         \regs[22][11] , \regs[22][10] , \regs[22][9] , \regs[22][8] ,
         \regs[22][7] , \regs[22][6] , \regs[22][5] , \regs[22][4] ,
         \regs[22][3] , \regs[22][2] , \regs[22][1] , \regs[22][0] ,
         \regs[21][31] , \regs[21][30] , \regs[21][29] , \regs[21][28] ,
         \regs[21][27] , \regs[21][26] , \regs[21][25] , \regs[21][24] ,
         \regs[21][23] , \regs[21][22] , \regs[21][21] , \regs[21][20] ,
         \regs[21][19] , \regs[21][18] , \regs[21][17] , \regs[21][16] ,
         \regs[21][15] , \regs[21][14] , \regs[21][13] , \regs[21][12] ,
         \regs[21][11] , \regs[21][10] , \regs[21][9] , \regs[21][8] ,
         \regs[21][7] , \regs[21][6] , \regs[21][5] , \regs[21][4] ,
         \regs[21][3] , \regs[21][2] , \regs[21][1] , \regs[21][0] ,
         \regs[20][31] , \regs[20][30] , \regs[20][29] , \regs[20][28] ,
         \regs[20][27] , \regs[20][26] , \regs[20][25] , \regs[20][24] ,
         \regs[20][23] , \regs[20][22] , \regs[20][21] , \regs[20][20] ,
         \regs[20][19] , \regs[20][18] , \regs[20][17] , \regs[20][16] ,
         \regs[20][15] , \regs[20][14] , \regs[20][13] , \regs[20][12] ,
         \regs[20][11] , \regs[20][10] , \regs[20][9] , \regs[20][8] ,
         \regs[20][7] , \regs[20][6] , \regs[20][5] , \regs[20][4] ,
         \regs[20][3] , \regs[20][2] , \regs[20][1] , \regs[20][0] ,
         \regs[19][31] , \regs[19][30] , \regs[19][29] , \regs[19][28] ,
         \regs[19][27] , \regs[19][26] , \regs[19][25] , \regs[19][24] ,
         \regs[19][23] , \regs[19][22] , \regs[19][21] , \regs[19][20] ,
         \regs[19][19] , \regs[19][18] , \regs[19][17] , \regs[19][16] ,
         \regs[19][15] , \regs[19][14] , \regs[19][13] , \regs[19][12] ,
         \regs[19][11] , \regs[19][10] , \regs[19][9] , \regs[19][8] ,
         \regs[19][7] , \regs[19][6] , \regs[19][5] , \regs[19][4] ,
         \regs[19][3] , \regs[19][2] , \regs[19][1] , \regs[19][0] ,
         \regs[18][31] , \regs[18][30] , \regs[18][29] , \regs[18][28] ,
         \regs[18][27] , \regs[18][26] , \regs[18][25] , \regs[18][24] ,
         \regs[18][23] , \regs[18][22] , \regs[18][21] , \regs[18][20] ,
         \regs[18][19] , \regs[18][18] , \regs[18][17] , \regs[18][16] ,
         \regs[18][15] , \regs[18][14] , \regs[18][13] , \regs[18][12] ,
         \regs[18][11] , \regs[18][10] , \regs[18][9] , \regs[18][8] ,
         \regs[18][7] , \regs[18][6] , \regs[18][5] , \regs[18][4] ,
         \regs[18][3] , \regs[18][2] , \regs[18][1] , \regs[18][0] ,
         \regs[17][31] , \regs[17][30] , \regs[17][29] , \regs[17][28] ,
         \regs[17][27] , \regs[17][26] , \regs[17][25] , \regs[17][24] ,
         \regs[17][23] , \regs[17][22] , \regs[17][21] , \regs[17][20] ,
         \regs[17][19] , \regs[17][18] , \regs[17][17] , \regs[17][16] ,
         \regs[17][15] , \regs[17][14] , \regs[17][13] , \regs[17][12] ,
         \regs[17][11] , \regs[17][10] , \regs[17][9] , \regs[17][8] ,
         \regs[17][7] , \regs[17][6] , \regs[17][5] , \regs[17][4] ,
         \regs[17][3] , \regs[17][2] , \regs[17][1] , \regs[17][0] ,
         \regs[16][31] , \regs[16][30] , \regs[16][29] , \regs[16][28] ,
         \regs[16][27] , \regs[16][26] , \regs[16][25] , \regs[16][24] ,
         \regs[16][23] , \regs[16][22] , \regs[16][21] , \regs[16][20] ,
         \regs[16][19] , \regs[16][18] , \regs[16][17] , \regs[16][16] ,
         \regs[16][15] , \regs[16][14] , \regs[16][13] , \regs[16][12] ,
         \regs[16][11] , \regs[16][10] , \regs[16][9] , \regs[16][8] ,
         \regs[16][7] , \regs[16][6] , \regs[16][5] , \regs[16][4] ,
         \regs[16][3] , \regs[16][2] , \regs[16][1] , \regs[16][0] ,
         \regs[15][31] , \regs[15][30] , \regs[15][29] , \regs[15][28] ,
         \regs[15][27] , \regs[15][26] , \regs[15][25] , \regs[15][24] ,
         \regs[15][23] , \regs[15][22] , \regs[15][21] , \regs[15][20] ,
         \regs[15][19] , \regs[15][18] , \regs[15][17] , \regs[15][16] ,
         \regs[15][15] , \regs[15][14] , \regs[15][13] , \regs[15][12] ,
         \regs[15][11] , \regs[15][10] , \regs[15][9] , \regs[15][8] ,
         \regs[15][7] , \regs[15][6] , \regs[15][5] , \regs[15][4] ,
         \regs[15][3] , \regs[15][2] , \regs[15][1] , \regs[15][0] ,
         \regs[14][31] , \regs[14][30] , \regs[14][29] , \regs[14][28] ,
         \regs[14][27] , \regs[14][26] , \regs[14][25] , \regs[14][24] ,
         \regs[14][23] , \regs[14][22] , \regs[14][21] , \regs[14][20] ,
         \regs[14][19] , \regs[14][18] , \regs[14][17] , \regs[14][16] ,
         \regs[14][15] , \regs[14][14] , \regs[14][13] , \regs[14][12] ,
         \regs[14][11] , \regs[14][10] , \regs[14][9] , \regs[14][8] ,
         \regs[14][7] , \regs[14][6] , \regs[14][5] , \regs[14][4] ,
         \regs[14][3] , \regs[14][2] , \regs[14][1] , \regs[14][0] ,
         \regs[13][31] , \regs[13][30] , \regs[13][29] , \regs[13][28] ,
         \regs[13][27] , \regs[13][26] , \regs[13][25] , \regs[13][24] ,
         \regs[13][23] , \regs[13][22] , \regs[13][21] , \regs[13][20] ,
         \regs[13][19] , \regs[13][18] , \regs[13][17] , \regs[13][16] ,
         \regs[13][15] , \regs[13][14] , \regs[13][13] , \regs[13][12] ,
         \regs[13][11] , \regs[13][10] , \regs[13][9] , \regs[13][8] ,
         \regs[13][7] , \regs[13][6] , \regs[13][5] , \regs[13][4] ,
         \regs[13][3] , \regs[13][2] , \regs[13][1] , \regs[13][0] ,
         \regs[12][31] , \regs[12][30] , \regs[12][29] , \regs[12][28] ,
         \regs[12][27] , \regs[12][26] , \regs[12][25] , \regs[12][24] ,
         \regs[12][23] , \regs[12][22] , \regs[12][21] , \regs[12][20] ,
         \regs[12][19] , \regs[12][18] , \regs[12][17] , \regs[12][16] ,
         \regs[12][15] , \regs[12][14] , \regs[12][13] , \regs[12][12] ,
         \regs[12][11] , \regs[12][10] , \regs[12][9] , \regs[12][8] ,
         \regs[12][7] , \regs[12][6] , \regs[12][5] , \regs[12][4] ,
         \regs[12][3] , \regs[12][2] , \regs[12][1] , \regs[12][0] ,
         \regs[11][31] , \regs[11][30] , \regs[11][29] , \regs[11][28] ,
         \regs[11][27] , \regs[11][26] , \regs[11][25] , \regs[11][24] ,
         \regs[11][23] , \regs[11][22] , \regs[11][21] , \regs[11][20] ,
         \regs[11][19] , \regs[11][18] , \regs[11][17] , \regs[11][16] ,
         \regs[11][15] , \regs[11][14] , \regs[11][13] , \regs[11][12] ,
         \regs[11][11] , \regs[11][10] , \regs[11][9] , \regs[11][8] ,
         \regs[11][7] , \regs[11][6] , \regs[11][5] , \regs[11][4] ,
         \regs[11][3] , \regs[11][2] , \regs[11][1] , \regs[11][0] ,
         \regs[10][31] , \regs[10][30] , \regs[10][29] , \regs[10][28] ,
         \regs[10][27] , \regs[10][26] , \regs[10][25] , \regs[10][24] ,
         \regs[10][23] , \regs[10][22] , \regs[10][21] , \regs[10][20] ,
         \regs[10][19] , \regs[10][18] , \regs[10][17] , \regs[10][16] ,
         \regs[10][15] , \regs[10][14] , \regs[10][13] , \regs[10][12] ,
         \regs[10][11] , \regs[10][10] , \regs[10][9] , \regs[10][8] ,
         \regs[10][7] , \regs[10][6] , \regs[10][5] , \regs[10][4] ,
         \regs[10][3] , \regs[10][2] , \regs[10][1] , \regs[10][0] ,
         \regs[9][31] , \regs[9][30] , \regs[9][29] , \regs[9][28] ,
         \regs[9][27] , \regs[9][26] , \regs[9][25] , \regs[9][24] ,
         \regs[9][23] , \regs[9][22] , \regs[9][21] , \regs[9][20] ,
         \regs[9][19] , \regs[9][18] , \regs[9][17] , \regs[9][16] ,
         \regs[9][15] , \regs[9][14] , \regs[9][13] , \regs[9][12] ,
         \regs[9][11] , \regs[9][10] , \regs[9][9] , \regs[9][8] ,
         \regs[9][7] , \regs[9][6] , \regs[9][5] , \regs[9][4] , \regs[9][3] ,
         \regs[9][2] , \regs[9][1] , \regs[9][0] , \regs[8][31] ,
         \regs[8][30] , \regs[8][29] , \regs[8][28] , \regs[8][27] ,
         \regs[8][26] , \regs[8][25] , \regs[8][24] , \regs[8][23] ,
         \regs[8][22] , \regs[8][21] , \regs[8][20] , \regs[8][19] ,
         \regs[8][18] , \regs[8][17] , \regs[8][16] , \regs[8][15] ,
         \regs[8][14] , \regs[8][13] , \regs[8][12] , \regs[8][11] ,
         \regs[8][10] , \regs[8][9] , \regs[8][8] , \regs[8][7] , \regs[8][6] ,
         \regs[8][5] , \regs[8][4] , \regs[8][3] , \regs[8][2] , \regs[8][1] ,
         \regs[8][0] , \regs[7][31] , \regs[7][30] , \regs[7][29] ,
         \regs[7][28] , \regs[7][27] , \regs[7][26] , \regs[7][25] ,
         \regs[7][24] , \regs[7][23] , \regs[7][22] , \regs[7][21] ,
         \regs[7][20] , \regs[7][19] , \regs[7][18] , \regs[7][17] ,
         \regs[7][16] , \regs[7][15] , \regs[7][14] , \regs[7][13] ,
         \regs[7][12] , \regs[7][11] , \regs[7][10] , \regs[7][9] ,
         \regs[7][8] , \regs[7][7] , \regs[7][6] , \regs[7][5] , \regs[7][4] ,
         \regs[7][3] , \regs[7][2] , \regs[7][1] , \regs[7][0] , \regs[6][31] ,
         \regs[6][30] , \regs[6][29] , \regs[6][28] , \regs[6][27] ,
         \regs[6][26] , \regs[6][25] , \regs[6][24] , \regs[6][23] ,
         \regs[6][22] , \regs[6][21] , \regs[6][20] , \regs[6][19] ,
         \regs[6][18] , \regs[6][17] , \regs[6][16] , \regs[6][15] ,
         \regs[6][14] , \regs[6][13] , \regs[6][12] , \regs[6][11] ,
         \regs[6][10] , \regs[6][9] , \regs[6][8] , \regs[6][7] , \regs[6][6] ,
         \regs[6][5] , \regs[6][4] , \regs[6][3] , \regs[6][2] , \regs[6][1] ,
         \regs[6][0] , \regs[5][31] , \regs[5][30] , \regs[5][29] ,
         \regs[5][28] , \regs[5][27] , \regs[5][26] , \regs[5][25] ,
         \regs[5][24] , \regs[5][23] , \regs[5][22] , \regs[5][21] ,
         \regs[5][20] , \regs[5][19] , \regs[5][18] , \regs[5][17] ,
         \regs[5][16] , \regs[5][15] , \regs[5][14] , \regs[5][13] ,
         \regs[5][12] , \regs[5][11] , \regs[5][10] , \regs[5][9] ,
         \regs[5][8] , \regs[5][7] , \regs[5][6] , \regs[5][5] , \regs[5][4] ,
         \regs[5][3] , \regs[5][2] , \regs[5][1] , \regs[5][0] , \regs[4][31] ,
         \regs[4][30] , \regs[4][29] , \regs[4][28] , \regs[4][27] ,
         \regs[4][26] , \regs[4][25] , \regs[4][24] , \regs[4][23] ,
         \regs[4][22] , \regs[4][21] , \regs[4][20] , \regs[4][19] ,
         \regs[4][18] , \regs[4][17] , \regs[4][16] , \regs[4][15] ,
         \regs[4][14] , \regs[4][13] , \regs[4][12] , \regs[4][11] ,
         \regs[4][10] , \regs[4][9] , \regs[4][8] , \regs[4][7] , \regs[4][6] ,
         \regs[4][5] , \regs[4][4] , \regs[4][3] , \regs[4][2] , \regs[4][1] ,
         \regs[4][0] , \regs[3][31] , \regs[3][30] , \regs[3][29] ,
         \regs[3][28] , \regs[3][27] , \regs[3][26] , \regs[3][25] ,
         \regs[3][24] , \regs[3][23] , \regs[3][22] , \regs[3][21] ,
         \regs[3][20] , \regs[3][19] , \regs[3][18] , \regs[3][17] ,
         \regs[3][16] , \regs[3][15] , \regs[3][14] , \regs[3][13] ,
         \regs[3][12] , \regs[3][11] , \regs[3][10] , \regs[3][9] ,
         \regs[3][8] , \regs[3][7] , \regs[3][6] , \regs[3][5] , \regs[3][4] ,
         \regs[3][3] , \regs[3][2] , \regs[3][1] , \regs[3][0] , \regs[2][31] ,
         \regs[2][30] , \regs[2][29] , \regs[2][28] , \regs[2][27] ,
         \regs[2][26] , \regs[2][25] , \regs[2][24] , \regs[2][23] ,
         \regs[2][22] , \regs[2][21] , \regs[2][20] , \regs[2][19] ,
         \regs[2][18] , \regs[2][17] , \regs[2][16] , \regs[2][15] ,
         \regs[2][14] , \regs[2][13] , \regs[2][12] , \regs[2][11] ,
         \regs[2][10] , \regs[2][9] , \regs[2][8] , \regs[2][7] , \regs[2][6] ,
         \regs[2][5] , \regs[2][4] , \regs[2][3] , \regs[2][2] , \regs[2][1] ,
         \regs[2][0] , \regs[1][31] , \regs[1][30] , \regs[1][29] ,
         \regs[1][28] , \regs[1][27] , \regs[1][26] , \regs[1][25] ,
         \regs[1][24] , \regs[1][23] , \regs[1][22] , \regs[1][21] ,
         \regs[1][20] , \regs[1][19] , \regs[1][18] , \regs[1][17] ,
         \regs[1][16] , \regs[1][15] , \regs[1][14] , \regs[1][13] ,
         \regs[1][12] , \regs[1][11] , \regs[1][10] , \regs[1][9] ,
         \regs[1][8] , \regs[1][7] , \regs[1][6] , \regs[1][5] , \regs[1][4] ,
         \regs[1][3] , \regs[1][2] , \regs[1][1] , \regs[1][0] , \regs[0][31] ,
         \regs[0][30] , \regs[0][29] , \regs[0][28] , \regs[0][27] ,
         \regs[0][26] , \regs[0][25] , \regs[0][24] , \regs[0][23] ,
         \regs[0][22] , \regs[0][21] , \regs[0][20] , \regs[0][19] ,
         \regs[0][18] , \regs[0][17] , \regs[0][16] , \regs[0][15] ,
         \regs[0][14] , \regs[0][13] , \regs[0][12] , \regs[0][11] ,
         \regs[0][10] , \regs[0][9] , \regs[0][8] , \regs[0][7] , \regs[0][6] ,
         \regs[0][5] , \regs[0][4] , \regs[0][3] , \regs[0][2] , \regs[0][1] ,
         \regs[0][0] , N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093,
         N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103,
         N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113,
         N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133,
         N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153,
         N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163,
         N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173,
         N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, n2, n6, n7,
         n8, n9, n10, n11, n12, n34, n35, n36, n38, n40, n42, n43, n44, n46,
         n50, n52, n56, n58, n61, n62, n64, n66, n67, n68, n70, n74, n76, n81,
         n83, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1, n3, n4,
         n5, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n37, n39, n41, n45, n47, n48,
         n49, n51, n53, n54, n55, n57, n59, n60, n63, n65, n69, n71, n72, n73,
         n75, n77, n78, n79, n80, n82, n84, n85, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227;
  assign N12 = addr1[0];
  assign N13 = addr1[1];
  assign N14 = addr1[2];
  assign N15 = addr1[3];
  assign N16 = addr1[4];
  assign N17 = addr2[0];
  assign N18 = addr2[1];
  assign N19 = addr2[2];
  assign N20 = addr2[3];
  assign N21 = addr2[4];
  assign N22 = addr_dst[0];
  assign N23 = addr_dst[1];
  assign N24 = addr_dst[2];
  assign N25 = addr_dst[3];
  assign N26 = addr_dst[4];

  DFFRHQX1 \regs_reg[29][31]  ( .D(n1045), .CK(clk), .RN(rst), .Q(
        \regs[29][31] ) );
  DFFRHQX1 \regs_reg[29][30]  ( .D(n1044), .CK(clk), .RN(rst), .Q(
        \regs[29][30] ) );
  DFFRHQX1 \regs_reg[29][29]  ( .D(n1043), .CK(clk), .RN(rst), .Q(
        \regs[29][29] ) );
  DFFRHQX1 \regs_reg[29][28]  ( .D(n1042), .CK(clk), .RN(rst), .Q(
        \regs[29][28] ) );
  DFFRHQX1 \regs_reg[29][27]  ( .D(n1041), .CK(clk), .RN(rst), .Q(
        \regs[29][27] ) );
  DFFRHQX1 \regs_reg[29][26]  ( .D(n1040), .CK(clk), .RN(rst), .Q(
        \regs[29][26] ) );
  DFFRHQX1 \regs_reg[29][25]  ( .D(n1039), .CK(clk), .RN(rst), .Q(
        \regs[29][25] ) );
  DFFRHQX1 \regs_reg[29][24]  ( .D(n1038), .CK(clk), .RN(rst), .Q(
        \regs[29][24] ) );
  DFFRHQX1 \regs_reg[29][15]  ( .D(n1029), .CK(clk), .RN(rst), .Q(
        \regs[29][15] ) );
  DFFRHQX1 \regs_reg[29][14]  ( .D(n1028), .CK(clk), .RN(rst), .Q(
        \regs[29][14] ) );
  DFFRHQX1 \regs_reg[29][13]  ( .D(n1027), .CK(clk), .RN(rst), .Q(
        \regs[29][13] ) );
  DFFRHQX1 \regs_reg[29][12]  ( .D(n1026), .CK(clk), .RN(rst), .Q(
        \regs[29][12] ) );
  DFFRHQX1 \regs_reg[29][11]  ( .D(n1025), .CK(clk), .RN(rst), .Q(
        \regs[29][11] ) );
  DFFRHQX1 \regs_reg[29][10]  ( .D(n1024), .CK(clk), .RN(rst), .Q(
        \regs[29][10] ) );
  DFFRHQX1 \regs_reg[29][9]  ( .D(n1023), .CK(clk), .RN(rst), .Q(\regs[29][9] ) );
  DFFRHQX1 \regs_reg[29][8]  ( .D(n1022), .CK(clk), .RN(rst), .Q(\regs[29][8] ) );
  DFFRHQX1 \regs_reg[29][7]  ( .D(n1021), .CK(clk), .RN(rst), .Q(\regs[29][7] ) );
  DFFRHQX1 \regs_reg[29][6]  ( .D(n1020), .CK(clk), .RN(rst), .Q(\regs[29][6] ) );
  DFFRHQX1 \regs_reg[29][5]  ( .D(n1019), .CK(clk), .RN(rst), .Q(\regs[29][5] ) );
  DFFRHQX1 \regs_reg[29][4]  ( .D(n1018), .CK(clk), .RN(rst), .Q(\regs[29][4] ) );
  DFFRHQX1 \regs_reg[29][3]  ( .D(n1017), .CK(clk), .RN(rst), .Q(\regs[29][3] ) );
  DFFRHQX1 \regs_reg[29][2]  ( .D(n1016), .CK(clk), .RN(rst), .Q(\regs[29][2] ) );
  DFFRHQX1 \regs_reg[29][1]  ( .D(n1015), .CK(clk), .RN(rst), .Q(\regs[29][1] ) );
  DFFRHQX1 \regs_reg[29][0]  ( .D(n1014), .CK(clk), .RN(rst), .Q(\regs[29][0] ) );
  DFFRHQX1 \regs_reg[25][31]  ( .D(n917), .CK(clk), .RN(rst), .Q(
        \regs[25][31] ) );
  DFFRHQX1 \regs_reg[25][30]  ( .D(n916), .CK(clk), .RN(rst), .Q(
        \regs[25][30] ) );
  DFFRHQX1 \regs_reg[25][29]  ( .D(n915), .CK(clk), .RN(rst), .Q(
        \regs[25][29] ) );
  DFFRHQX1 \regs_reg[25][28]  ( .D(n914), .CK(clk), .RN(rst), .Q(
        \regs[25][28] ) );
  DFFRHQX1 \regs_reg[25][27]  ( .D(n913), .CK(clk), .RN(rst), .Q(
        \regs[25][27] ) );
  DFFRHQX1 \regs_reg[25][26]  ( .D(n912), .CK(clk), .RN(rst), .Q(
        \regs[25][26] ) );
  DFFRHQX1 \regs_reg[25][25]  ( .D(n911), .CK(clk), .RN(rst), .Q(
        \regs[25][25] ) );
  DFFRHQX1 \regs_reg[25][24]  ( .D(n910), .CK(clk), .RN(rst), .Q(
        \regs[25][24] ) );
  DFFRHQX1 \regs_reg[25][15]  ( .D(n901), .CK(clk), .RN(rst), .Q(
        \regs[25][15] ) );
  DFFRHQX1 \regs_reg[25][14]  ( .D(n900), .CK(clk), .RN(rst), .Q(
        \regs[25][14] ) );
  DFFRHQX1 \regs_reg[25][13]  ( .D(n899), .CK(clk), .RN(rst), .Q(
        \regs[25][13] ) );
  DFFRHQX1 \regs_reg[25][12]  ( .D(n898), .CK(clk), .RN(rst), .Q(
        \regs[25][12] ) );
  DFFRHQX1 \regs_reg[25][11]  ( .D(n897), .CK(clk), .RN(rst), .Q(
        \regs[25][11] ) );
  DFFRHQX1 \regs_reg[25][10]  ( .D(n896), .CK(clk), .RN(rst), .Q(
        \regs[25][10] ) );
  DFFRHQX1 \regs_reg[25][9]  ( .D(n895), .CK(clk), .RN(rst), .Q(\regs[25][9] )
         );
  DFFRHQX1 \regs_reg[25][8]  ( .D(n894), .CK(clk), .RN(rst), .Q(\regs[25][8] )
         );
  DFFRHQX1 \regs_reg[25][7]  ( .D(n893), .CK(clk), .RN(rst), .Q(\regs[25][7] )
         );
  DFFRHQX1 \regs_reg[25][6]  ( .D(n892), .CK(clk), .RN(rst), .Q(\regs[25][6] )
         );
  DFFRHQX1 \regs_reg[25][5]  ( .D(n891), .CK(clk), .RN(rst), .Q(\regs[25][5] )
         );
  DFFRHQX1 \regs_reg[25][4]  ( .D(n890), .CK(clk), .RN(rst), .Q(\regs[25][4] )
         );
  DFFRHQX1 \regs_reg[25][3]  ( .D(n889), .CK(clk), .RN(rst), .Q(\regs[25][3] )
         );
  DFFRHQX1 \regs_reg[25][2]  ( .D(n888), .CK(clk), .RN(rst), .Q(\regs[25][2] )
         );
  DFFRHQX1 \regs_reg[25][1]  ( .D(n887), .CK(clk), .RN(rst), .Q(\regs[25][1] )
         );
  DFFRHQX1 \regs_reg[25][0]  ( .D(n886), .CK(clk), .RN(rst), .Q(\regs[25][0] )
         );
  DFFRHQX1 \regs_reg[21][31]  ( .D(n789), .CK(clk), .RN(rst), .Q(
        \regs[21][31] ) );
  DFFRHQX1 \regs_reg[21][30]  ( .D(n788), .CK(clk), .RN(rst), .Q(
        \regs[21][30] ) );
  DFFRHQX1 \regs_reg[21][29]  ( .D(n787), .CK(clk), .RN(rst), .Q(
        \regs[21][29] ) );
  DFFRHQX1 \regs_reg[21][28]  ( .D(n786), .CK(clk), .RN(rst), .Q(
        \regs[21][28] ) );
  DFFRHQX1 \regs_reg[21][27]  ( .D(n785), .CK(clk), .RN(rst), .Q(
        \regs[21][27] ) );
  DFFRHQX1 \regs_reg[21][26]  ( .D(n784), .CK(clk), .RN(rst), .Q(
        \regs[21][26] ) );
  DFFRHQX1 \regs_reg[21][25]  ( .D(n783), .CK(clk), .RN(rst), .Q(
        \regs[21][25] ) );
  DFFRHQX1 \regs_reg[21][24]  ( .D(n782), .CK(clk), .RN(rst), .Q(
        \regs[21][24] ) );
  DFFRHQX1 \regs_reg[21][15]  ( .D(n773), .CK(clk), .RN(rst), .Q(
        \regs[21][15] ) );
  DFFRHQX1 \regs_reg[21][14]  ( .D(n772), .CK(clk), .RN(rst), .Q(
        \regs[21][14] ) );
  DFFRHQX1 \regs_reg[21][13]  ( .D(n771), .CK(clk), .RN(rst), .Q(
        \regs[21][13] ) );
  DFFRHQX1 \regs_reg[21][12]  ( .D(n770), .CK(clk), .RN(rst), .Q(
        \regs[21][12] ) );
  DFFRHQX1 \regs_reg[21][11]  ( .D(n769), .CK(clk), .RN(rst), .Q(
        \regs[21][11] ) );
  DFFRHQX1 \regs_reg[21][10]  ( .D(n768), .CK(clk), .RN(rst), .Q(
        \regs[21][10] ) );
  DFFRHQX1 \regs_reg[21][9]  ( .D(n767), .CK(clk), .RN(rst), .Q(\regs[21][9] )
         );
  DFFRHQX1 \regs_reg[21][8]  ( .D(n766), .CK(clk), .RN(rst), .Q(\regs[21][8] )
         );
  DFFRHQX1 \regs_reg[21][7]  ( .D(n765), .CK(clk), .RN(rst), .Q(\regs[21][7] )
         );
  DFFRHQX1 \regs_reg[21][6]  ( .D(n764), .CK(clk), .RN(rst), .Q(\regs[21][6] )
         );
  DFFRHQX1 \regs_reg[21][5]  ( .D(n763), .CK(clk), .RN(rst), .Q(\regs[21][5] )
         );
  DFFRHQX1 \regs_reg[21][4]  ( .D(n762), .CK(clk), .RN(rst), .Q(\regs[21][4] )
         );
  DFFRHQX1 \regs_reg[21][3]  ( .D(n761), .CK(clk), .RN(rst), .Q(\regs[21][3] )
         );
  DFFRHQX1 \regs_reg[21][2]  ( .D(n760), .CK(clk), .RN(rst), .Q(\regs[21][2] )
         );
  DFFRHQX1 \regs_reg[21][1]  ( .D(n759), .CK(clk), .RN(rst), .Q(\regs[21][1] )
         );
  DFFRHQX1 \regs_reg[21][0]  ( .D(n758), .CK(clk), .RN(rst), .Q(\regs[21][0] )
         );
  DFFRHQX1 \regs_reg[17][31]  ( .D(n661), .CK(clk), .RN(rst), .Q(
        \regs[17][31] ) );
  DFFRHQX1 \regs_reg[17][30]  ( .D(n660), .CK(clk), .RN(rst), .Q(
        \regs[17][30] ) );
  DFFRHQX1 \regs_reg[17][29]  ( .D(n659), .CK(clk), .RN(rst), .Q(
        \regs[17][29] ) );
  DFFRHQX1 \regs_reg[17][28]  ( .D(n658), .CK(clk), .RN(rst), .Q(
        \regs[17][28] ) );
  DFFRHQX1 \regs_reg[17][27]  ( .D(n657), .CK(clk), .RN(rst), .Q(
        \regs[17][27] ) );
  DFFRHQX1 \regs_reg[17][26]  ( .D(n656), .CK(clk), .RN(rst), .Q(
        \regs[17][26] ) );
  DFFRHQX1 \regs_reg[17][25]  ( .D(n655), .CK(clk), .RN(rst), .Q(
        \regs[17][25] ) );
  DFFRHQX1 \regs_reg[17][24]  ( .D(n654), .CK(clk), .RN(rst), .Q(
        \regs[17][24] ) );
  DFFRHQX1 \regs_reg[17][19]  ( .D(n649), .CK(clk), .RN(rst), .Q(
        \regs[17][19] ) );
  DFFRHQX1 \regs_reg[17][15]  ( .D(n645), .CK(clk), .RN(rst), .Q(
        \regs[17][15] ) );
  DFFRHQX1 \regs_reg[17][14]  ( .D(n644), .CK(clk), .RN(rst), .Q(
        \regs[17][14] ) );
  DFFRHQX1 \regs_reg[17][13]  ( .D(n643), .CK(clk), .RN(rst), .Q(
        \regs[17][13] ) );
  DFFRHQX1 \regs_reg[17][12]  ( .D(n642), .CK(clk), .RN(rst), .Q(
        \regs[17][12] ) );
  DFFRHQX1 \regs_reg[17][11]  ( .D(n641), .CK(clk), .RN(rst), .Q(
        \regs[17][11] ) );
  DFFRHQX1 \regs_reg[17][10]  ( .D(n640), .CK(clk), .RN(rst), .Q(
        \regs[17][10] ) );
  DFFRHQX1 \regs_reg[17][9]  ( .D(n639), .CK(clk), .RN(rst), .Q(\regs[17][9] )
         );
  DFFRHQX1 \regs_reg[17][8]  ( .D(n638), .CK(clk), .RN(rst), .Q(\regs[17][8] )
         );
  DFFRHQX1 \regs_reg[17][7]  ( .D(n637), .CK(clk), .RN(rst), .Q(\regs[17][7] )
         );
  DFFRHQX1 \regs_reg[17][6]  ( .D(n636), .CK(clk), .RN(rst), .Q(\regs[17][6] )
         );
  DFFRHQX1 \regs_reg[17][5]  ( .D(n635), .CK(clk), .RN(rst), .Q(\regs[17][5] )
         );
  DFFRHQX1 \regs_reg[17][4]  ( .D(n634), .CK(clk), .RN(rst), .Q(\regs[17][4] )
         );
  DFFRHQX1 \regs_reg[17][3]  ( .D(n633), .CK(clk), .RN(rst), .Q(\regs[17][3] )
         );
  DFFRHQX1 \regs_reg[17][2]  ( .D(n632), .CK(clk), .RN(rst), .Q(\regs[17][2] )
         );
  DFFRHQX1 \regs_reg[17][1]  ( .D(n631), .CK(clk), .RN(rst), .Q(\regs[17][1] )
         );
  DFFRHQX1 \regs_reg[17][0]  ( .D(n630), .CK(clk), .RN(rst), .Q(\regs[17][0] )
         );
  DFFRHQX1 \regs_reg[13][31]  ( .D(n533), .CK(clk), .RN(rst), .Q(
        \regs[13][31] ) );
  DFFRHQX1 \regs_reg[13][30]  ( .D(n532), .CK(clk), .RN(rst), .Q(
        \regs[13][30] ) );
  DFFRHQX1 \regs_reg[13][29]  ( .D(n531), .CK(clk), .RN(rst), .Q(
        \regs[13][29] ) );
  DFFRHQX1 \regs_reg[13][28]  ( .D(n530), .CK(clk), .RN(rst), .Q(
        \regs[13][28] ) );
  DFFRHQX1 \regs_reg[13][27]  ( .D(n529), .CK(clk), .RN(rst), .Q(
        \regs[13][27] ) );
  DFFRHQX1 \regs_reg[13][26]  ( .D(n528), .CK(clk), .RN(rst), .Q(
        \regs[13][26] ) );
  DFFRHQX1 \regs_reg[13][25]  ( .D(n527), .CK(clk), .RN(rst), .Q(
        \regs[13][25] ) );
  DFFRHQX1 \regs_reg[13][24]  ( .D(n526), .CK(clk), .RN(rst), .Q(
        \regs[13][24] ) );
  DFFRHQX1 \regs_reg[13][15]  ( .D(n517), .CK(clk), .RN(rst), .Q(
        \regs[13][15] ) );
  DFFRHQX1 \regs_reg[13][14]  ( .D(n516), .CK(clk), .RN(rst), .Q(
        \regs[13][14] ) );
  DFFRHQX1 \regs_reg[13][13]  ( .D(n515), .CK(clk), .RN(rst), .Q(
        \regs[13][13] ) );
  DFFRHQX1 \regs_reg[13][12]  ( .D(n514), .CK(clk), .RN(rst), .Q(
        \regs[13][12] ) );
  DFFRHQX1 \regs_reg[13][11]  ( .D(n513), .CK(clk), .RN(rst), .Q(
        \regs[13][11] ) );
  DFFRHQX1 \regs_reg[13][10]  ( .D(n512), .CK(clk), .RN(rst), .Q(
        \regs[13][10] ) );
  DFFRHQX1 \regs_reg[13][9]  ( .D(n511), .CK(clk), .RN(rst), .Q(\regs[13][9] )
         );
  DFFRHQX1 \regs_reg[13][8]  ( .D(n510), .CK(clk), .RN(rst), .Q(\regs[13][8] )
         );
  DFFRHQX1 \regs_reg[13][7]  ( .D(n509), .CK(clk), .RN(rst), .Q(\regs[13][7] )
         );
  DFFRHQX1 \regs_reg[13][6]  ( .D(n508), .CK(clk), .RN(rst), .Q(\regs[13][6] )
         );
  DFFRHQX1 \regs_reg[13][5]  ( .D(n507), .CK(clk), .RN(rst), .Q(\regs[13][5] )
         );
  DFFRHQX1 \regs_reg[13][4]  ( .D(n506), .CK(clk), .RN(rst), .Q(\regs[13][4] )
         );
  DFFRHQX1 \regs_reg[13][3]  ( .D(n505), .CK(clk), .RN(rst), .Q(\regs[13][3] )
         );
  DFFRHQX1 \regs_reg[13][2]  ( .D(n504), .CK(clk), .RN(rst), .Q(\regs[13][2] )
         );
  DFFRHQX1 \regs_reg[13][1]  ( .D(n503), .CK(clk), .RN(rst), .Q(\regs[13][1] )
         );
  DFFRHQX1 \regs_reg[13][0]  ( .D(n502), .CK(clk), .RN(rst), .Q(\regs[13][0] )
         );
  DFFRHQX1 \regs_reg[9][31]  ( .D(n405), .CK(clk), .RN(rst), .Q(\regs[9][31] )
         );
  DFFRHQX1 \regs_reg[9][30]  ( .D(n404), .CK(clk), .RN(rst), .Q(\regs[9][30] )
         );
  DFFRHQX1 \regs_reg[9][29]  ( .D(n403), .CK(clk), .RN(rst), .Q(\regs[9][29] )
         );
  DFFRHQX1 \regs_reg[9][28]  ( .D(n402), .CK(clk), .RN(rst), .Q(\regs[9][28] )
         );
  DFFRHQX1 \regs_reg[9][27]  ( .D(n401), .CK(clk), .RN(rst), .Q(\regs[9][27] )
         );
  DFFRHQX1 \regs_reg[9][26]  ( .D(n400), .CK(clk), .RN(rst), .Q(\regs[9][26] )
         );
  DFFRHQX1 \regs_reg[9][25]  ( .D(n399), .CK(clk), .RN(rst), .Q(\regs[9][25] )
         );
  DFFRHQX1 \regs_reg[9][24]  ( .D(n398), .CK(clk), .RN(rst), .Q(\regs[9][24] )
         );
  DFFRHQX1 \regs_reg[9][19]  ( .D(n393), .CK(clk), .RN(rst), .Q(\regs[9][19] )
         );
  DFFRHQX1 \regs_reg[9][15]  ( .D(n389), .CK(clk), .RN(rst), .Q(\regs[9][15] )
         );
  DFFRHQX1 \regs_reg[9][14]  ( .D(n388), .CK(clk), .RN(rst), .Q(\regs[9][14] )
         );
  DFFRHQX1 \regs_reg[9][13]  ( .D(n387), .CK(clk), .RN(rst), .Q(\regs[9][13] )
         );
  DFFRHQX1 \regs_reg[9][12]  ( .D(n386), .CK(clk), .RN(rst), .Q(\regs[9][12] )
         );
  DFFRHQX1 \regs_reg[9][11]  ( .D(n385), .CK(clk), .RN(rst), .Q(\regs[9][11] )
         );
  DFFRHQX1 \regs_reg[9][10]  ( .D(n384), .CK(clk), .RN(rst), .Q(\regs[9][10] )
         );
  DFFRHQX1 \regs_reg[9][9]  ( .D(n383), .CK(clk), .RN(rst), .Q(\regs[9][9] )
         );
  DFFRHQX1 \regs_reg[9][8]  ( .D(n382), .CK(clk), .RN(rst), .Q(\regs[9][8] )
         );
  DFFRHQX1 \regs_reg[9][7]  ( .D(n381), .CK(clk), .RN(rst), .Q(\regs[9][7] )
         );
  DFFRHQX1 \regs_reg[9][6]  ( .D(n380), .CK(clk), .RN(rst), .Q(\regs[9][6] )
         );
  DFFRHQX1 \regs_reg[9][5]  ( .D(n379), .CK(clk), .RN(rst), .Q(\regs[9][5] )
         );
  DFFRHQX1 \regs_reg[9][4]  ( .D(n378), .CK(clk), .RN(rst), .Q(\regs[9][4] )
         );
  DFFRHQX1 \regs_reg[9][3]  ( .D(n377), .CK(clk), .RN(rst), .Q(\regs[9][3] )
         );
  DFFRHQX1 \regs_reg[9][2]  ( .D(n376), .CK(clk), .RN(rst), .Q(\regs[9][2] )
         );
  DFFRHQX1 \regs_reg[9][1]  ( .D(n375), .CK(clk), .RN(rst), .Q(\regs[9][1] )
         );
  DFFRHQX1 \regs_reg[9][0]  ( .D(n374), .CK(clk), .RN(rst), .Q(\regs[9][0] )
         );
  DFFRHQX1 \regs_reg[5][31]  ( .D(n277), .CK(clk), .RN(rst), .Q(\regs[5][31] )
         );
  DFFRHQX1 \regs_reg[5][30]  ( .D(n276), .CK(clk), .RN(rst), .Q(\regs[5][30] )
         );
  DFFRHQX1 \regs_reg[5][29]  ( .D(n275), .CK(clk), .RN(rst), .Q(\regs[5][29] )
         );
  DFFRHQX1 \regs_reg[5][28]  ( .D(n274), .CK(clk), .RN(rst), .Q(\regs[5][28] )
         );
  DFFRHQX1 \regs_reg[5][27]  ( .D(n273), .CK(clk), .RN(rst), .Q(\regs[5][27] )
         );
  DFFRHQX1 \regs_reg[5][26]  ( .D(n272), .CK(clk), .RN(rst), .Q(\regs[5][26] )
         );
  DFFRHQX1 \regs_reg[5][25]  ( .D(n271), .CK(clk), .RN(rst), .Q(\regs[5][25] )
         );
  DFFRHQX1 \regs_reg[5][24]  ( .D(n270), .CK(clk), .RN(rst), .Q(\regs[5][24] )
         );
  DFFRHQX1 \regs_reg[5][19]  ( .D(n265), .CK(clk), .RN(rst), .Q(\regs[5][19] )
         );
  DFFRHQX1 \regs_reg[5][15]  ( .D(n261), .CK(clk), .RN(rst), .Q(\regs[5][15] )
         );
  DFFRHQX1 \regs_reg[5][14]  ( .D(n260), .CK(clk), .RN(rst), .Q(\regs[5][14] )
         );
  DFFRHQX1 \regs_reg[5][13]  ( .D(n259), .CK(clk), .RN(rst), .Q(\regs[5][13] )
         );
  DFFRHQX1 \regs_reg[5][12]  ( .D(n258), .CK(clk), .RN(rst), .Q(\regs[5][12] )
         );
  DFFRHQX1 \regs_reg[5][11]  ( .D(n257), .CK(clk), .RN(rst), .Q(\regs[5][11] )
         );
  DFFRHQX1 \regs_reg[5][10]  ( .D(n256), .CK(clk), .RN(rst), .Q(\regs[5][10] )
         );
  DFFRHQX1 \regs_reg[5][9]  ( .D(n255), .CK(clk), .RN(rst), .Q(\regs[5][9] )
         );
  DFFRHQX1 \regs_reg[5][8]  ( .D(n254), .CK(clk), .RN(rst), .Q(\regs[5][8] )
         );
  DFFRHQX1 \regs_reg[5][7]  ( .D(n253), .CK(clk), .RN(rst), .Q(\regs[5][7] )
         );
  DFFRHQX1 \regs_reg[5][6]  ( .D(n252), .CK(clk), .RN(rst), .Q(\regs[5][6] )
         );
  DFFRHQX1 \regs_reg[5][5]  ( .D(n251), .CK(clk), .RN(rst), .Q(\regs[5][5] )
         );
  DFFRHQX1 \regs_reg[5][4]  ( .D(n250), .CK(clk), .RN(rst), .Q(\regs[5][4] )
         );
  DFFRHQX1 \regs_reg[5][3]  ( .D(n249), .CK(clk), .RN(rst), .Q(\regs[5][3] )
         );
  DFFRHQX1 \regs_reg[5][2]  ( .D(n248), .CK(clk), .RN(rst), .Q(\regs[5][2] )
         );
  DFFRHQX1 \regs_reg[5][1]  ( .D(n247), .CK(clk), .RN(rst), .Q(\regs[5][1] )
         );
  DFFRHQX1 \regs_reg[5][0]  ( .D(n246), .CK(clk), .RN(rst), .Q(\regs[5][0] )
         );
  DFFRHQX1 \regs_reg[1][31]  ( .D(n149), .CK(clk), .RN(rst), .Q(\regs[1][31] )
         );
  DFFRHQX1 \regs_reg[1][30]  ( .D(n148), .CK(clk), .RN(rst), .Q(\regs[1][30] )
         );
  DFFRHQX1 \regs_reg[1][29]  ( .D(n147), .CK(clk), .RN(rst), .Q(\regs[1][29] )
         );
  DFFRHQX1 \regs_reg[1][28]  ( .D(n146), .CK(clk), .RN(rst), .Q(\regs[1][28] )
         );
  DFFRHQX1 \regs_reg[1][27]  ( .D(n145), .CK(clk), .RN(rst), .Q(\regs[1][27] )
         );
  DFFRHQX1 \regs_reg[1][26]  ( .D(n144), .CK(clk), .RN(rst), .Q(\regs[1][26] )
         );
  DFFRHQX1 \regs_reg[1][25]  ( .D(n143), .CK(clk), .RN(rst), .Q(\regs[1][25] )
         );
  DFFRHQX1 \regs_reg[1][24]  ( .D(n142), .CK(clk), .RN(rst), .Q(\regs[1][24] )
         );
  DFFRHQX1 \regs_reg[1][19]  ( .D(n137), .CK(clk), .RN(rst), .Q(\regs[1][19] )
         );
  DFFRHQX1 \regs_reg[1][18]  ( .D(n136), .CK(clk), .RN(rst), .Q(\regs[1][18] )
         );
  DFFRHQX1 \regs_reg[1][15]  ( .D(n133), .CK(clk), .RN(rst), .Q(\regs[1][15] )
         );
  DFFRHQX1 \regs_reg[1][14]  ( .D(n132), .CK(clk), .RN(rst), .Q(\regs[1][14] )
         );
  DFFRHQX1 \regs_reg[1][13]  ( .D(n131), .CK(clk), .RN(rst), .Q(\regs[1][13] )
         );
  DFFRHQX1 \regs_reg[1][12]  ( .D(n130), .CK(clk), .RN(rst), .Q(\regs[1][12] )
         );
  DFFRHQX1 \regs_reg[1][11]  ( .D(n129), .CK(clk), .RN(rst), .Q(\regs[1][11] )
         );
  DFFRHQX1 \regs_reg[1][10]  ( .D(n128), .CK(clk), .RN(rst), .Q(\regs[1][10] )
         );
  DFFRHQX1 \regs_reg[1][9]  ( .D(n127), .CK(clk), .RN(rst), .Q(\regs[1][9] )
         );
  DFFRHQX1 \regs_reg[1][8]  ( .D(n126), .CK(clk), .RN(rst), .Q(\regs[1][8] )
         );
  DFFRHQX1 \regs_reg[1][7]  ( .D(n125), .CK(clk), .RN(rst), .Q(\regs[1][7] )
         );
  DFFRHQX1 \regs_reg[1][6]  ( .D(n124), .CK(clk), .RN(rst), .Q(\regs[1][6] )
         );
  DFFRHQX1 \regs_reg[1][5]  ( .D(n123), .CK(clk), .RN(rst), .Q(\regs[1][5] )
         );
  DFFRHQX1 \regs_reg[1][4]  ( .D(n122), .CK(clk), .RN(rst), .Q(\regs[1][4] )
         );
  DFFRHQX1 \regs_reg[1][3]  ( .D(n121), .CK(clk), .RN(rst), .Q(\regs[1][3] )
         );
  DFFRHQX1 \regs_reg[1][2]  ( .D(n120), .CK(clk), .RN(rst), .Q(\regs[1][2] )
         );
  DFFRHQX1 \regs_reg[1][1]  ( .D(n119), .CK(clk), .RN(rst), .Q(\regs[1][1] )
         );
  DFFRHQX1 \regs_reg[1][0]  ( .D(n118), .CK(clk), .RN(rst), .Q(\regs[1][0] )
         );
  DFFRHQX1 \regs_reg[31][31]  ( .D(n1109), .CK(clk), .RN(rst), .Q(
        \regs[31][31] ) );
  DFFRHQX1 \regs_reg[31][30]  ( .D(n1108), .CK(clk), .RN(rst), .Q(
        \regs[31][30] ) );
  DFFRHQX1 \regs_reg[31][29]  ( .D(n1107), .CK(clk), .RN(rst), .Q(
        \regs[31][29] ) );
  DFFRHQX1 \regs_reg[31][28]  ( .D(n1106), .CK(clk), .RN(rst), .Q(
        \regs[31][28] ) );
  DFFRHQX1 \regs_reg[31][27]  ( .D(n1105), .CK(clk), .RN(rst), .Q(
        \regs[31][27] ) );
  DFFRHQX1 \regs_reg[31][26]  ( .D(n1104), .CK(clk), .RN(rst), .Q(
        \regs[31][26] ) );
  DFFRHQX1 \regs_reg[31][25]  ( .D(n1103), .CK(clk), .RN(rst), .Q(
        \regs[31][25] ) );
  DFFRHQX1 \regs_reg[31][24]  ( .D(n1102), .CK(clk), .RN(rst), .Q(
        \regs[31][24] ) );
  DFFRHQX1 \regs_reg[31][15]  ( .D(n1093), .CK(clk), .RN(rst), .Q(
        \regs[31][15] ) );
  DFFRHQX1 \regs_reg[31][14]  ( .D(n1092), .CK(clk), .RN(rst), .Q(
        \regs[31][14] ) );
  DFFRHQX1 \regs_reg[31][13]  ( .D(n1091), .CK(clk), .RN(rst), .Q(
        \regs[31][13] ) );
  DFFRHQX1 \regs_reg[31][12]  ( .D(n1090), .CK(clk), .RN(rst), .Q(
        \regs[31][12] ) );
  DFFRHQX1 \regs_reg[31][11]  ( .D(n1089), .CK(clk), .RN(rst), .Q(
        \regs[31][11] ) );
  DFFRHQX1 \regs_reg[31][10]  ( .D(n1088), .CK(clk), .RN(rst), .Q(
        \regs[31][10] ) );
  DFFRHQX1 \regs_reg[31][9]  ( .D(n1087), .CK(clk), .RN(rst), .Q(\regs[31][9] ) );
  DFFRHQX1 \regs_reg[31][8]  ( .D(n1086), .CK(clk), .RN(rst), .Q(\regs[31][8] ) );
  DFFRHQX1 \regs_reg[31][7]  ( .D(n1085), .CK(clk), .RN(rst), .Q(\regs[31][7] ) );
  DFFRHQX1 \regs_reg[31][6]  ( .D(n1084), .CK(clk), .RN(rst), .Q(\regs[31][6] ) );
  DFFRHQX1 \regs_reg[31][5]  ( .D(n1083), .CK(clk), .RN(rst), .Q(\regs[31][5] ) );
  DFFRHQX1 \regs_reg[31][4]  ( .D(n1082), .CK(clk), .RN(rst), .Q(\regs[31][4] ) );
  DFFRHQX1 \regs_reg[31][3]  ( .D(n1081), .CK(clk), .RN(rst), .Q(\regs[31][3] ) );
  DFFRHQX1 \regs_reg[31][2]  ( .D(n1080), .CK(clk), .RN(rst), .Q(\regs[31][2] ) );
  DFFRHQX1 \regs_reg[31][1]  ( .D(n1079), .CK(clk), .RN(rst), .Q(\regs[31][1] ) );
  DFFRHQX1 \regs_reg[31][0]  ( .D(n1078), .CK(clk), .RN(rst), .Q(\regs[31][0] ) );
  DFFRHQX1 \regs_reg[27][31]  ( .D(n981), .CK(clk), .RN(rst), .Q(
        \regs[27][31] ) );
  DFFRHQX1 \regs_reg[27][30]  ( .D(n980), .CK(clk), .RN(rst), .Q(
        \regs[27][30] ) );
  DFFRHQX1 \regs_reg[27][29]  ( .D(n979), .CK(clk), .RN(rst), .Q(
        \regs[27][29] ) );
  DFFRHQX1 \regs_reg[27][28]  ( .D(n978), .CK(clk), .RN(rst), .Q(
        \regs[27][28] ) );
  DFFRHQX1 \regs_reg[27][27]  ( .D(n977), .CK(clk), .RN(rst), .Q(
        \regs[27][27] ) );
  DFFRHQX1 \regs_reg[27][26]  ( .D(n976), .CK(clk), .RN(rst), .Q(
        \regs[27][26] ) );
  DFFRHQX1 \regs_reg[27][25]  ( .D(n975), .CK(clk), .RN(rst), .Q(
        \regs[27][25] ) );
  DFFRHQX1 \regs_reg[27][24]  ( .D(n974), .CK(clk), .RN(rst), .Q(
        \regs[27][24] ) );
  DFFRHQX1 \regs_reg[27][15]  ( .D(n965), .CK(clk), .RN(rst), .Q(
        \regs[27][15] ) );
  DFFRHQX1 \regs_reg[27][14]  ( .D(n964), .CK(clk), .RN(rst), .Q(
        \regs[27][14] ) );
  DFFRHQX1 \regs_reg[27][13]  ( .D(n963), .CK(clk), .RN(rst), .Q(
        \regs[27][13] ) );
  DFFRHQX1 \regs_reg[27][12]  ( .D(n962), .CK(clk), .RN(rst), .Q(
        \regs[27][12] ) );
  DFFRHQX1 \regs_reg[27][11]  ( .D(n961), .CK(clk), .RN(rst), .Q(
        \regs[27][11] ) );
  DFFRHQX1 \regs_reg[27][10]  ( .D(n960), .CK(clk), .RN(rst), .Q(
        \regs[27][10] ) );
  DFFRHQX1 \regs_reg[27][9]  ( .D(n959), .CK(clk), .RN(rst), .Q(\regs[27][9] )
         );
  DFFRHQX1 \regs_reg[27][8]  ( .D(n958), .CK(clk), .RN(rst), .Q(\regs[27][8] )
         );
  DFFRHQX1 \regs_reg[27][7]  ( .D(n957), .CK(clk), .RN(rst), .Q(\regs[27][7] )
         );
  DFFRHQX1 \regs_reg[27][6]  ( .D(n956), .CK(clk), .RN(rst), .Q(\regs[27][6] )
         );
  DFFRHQX1 \regs_reg[27][5]  ( .D(n955), .CK(clk), .RN(rst), .Q(\regs[27][5] )
         );
  DFFRHQX1 \regs_reg[27][4]  ( .D(n954), .CK(clk), .RN(rst), .Q(\regs[27][4] )
         );
  DFFRHQX1 \regs_reg[27][3]  ( .D(n953), .CK(clk), .RN(rst), .Q(\regs[27][3] )
         );
  DFFRHQX1 \regs_reg[27][2]  ( .D(n952), .CK(clk), .RN(rst), .Q(\regs[27][2] )
         );
  DFFRHQX1 \regs_reg[27][1]  ( .D(n951), .CK(clk), .RN(rst), .Q(\regs[27][1] )
         );
  DFFRHQX1 \regs_reg[27][0]  ( .D(n950), .CK(clk), .RN(rst), .Q(\regs[27][0] )
         );
  DFFRHQX1 \regs_reg[23][31]  ( .D(n853), .CK(clk), .RN(rst), .Q(
        \regs[23][31] ) );
  DFFRHQX1 \regs_reg[23][30]  ( .D(n852), .CK(clk), .RN(rst), .Q(
        \regs[23][30] ) );
  DFFRHQX1 \regs_reg[23][29]  ( .D(n851), .CK(clk), .RN(rst), .Q(
        \regs[23][29] ) );
  DFFRHQX1 \regs_reg[23][28]  ( .D(n850), .CK(clk), .RN(rst), .Q(
        \regs[23][28] ) );
  DFFRHQX1 \regs_reg[23][27]  ( .D(n849), .CK(clk), .RN(rst), .Q(
        \regs[23][27] ) );
  DFFRHQX1 \regs_reg[23][26]  ( .D(n848), .CK(clk), .RN(rst), .Q(
        \regs[23][26] ) );
  DFFRHQX1 \regs_reg[23][25]  ( .D(n847), .CK(clk), .RN(rst), .Q(
        \regs[23][25] ) );
  DFFRHQX1 \regs_reg[23][24]  ( .D(n846), .CK(clk), .RN(rst), .Q(
        \regs[23][24] ) );
  DFFRHQX1 \regs_reg[23][15]  ( .D(n837), .CK(clk), .RN(rst), .Q(
        \regs[23][15] ) );
  DFFRHQX1 \regs_reg[23][14]  ( .D(n836), .CK(clk), .RN(rst), .Q(
        \regs[23][14] ) );
  DFFRHQX1 \regs_reg[23][13]  ( .D(n835), .CK(clk), .RN(rst), .Q(
        \regs[23][13] ) );
  DFFRHQX1 \regs_reg[23][12]  ( .D(n834), .CK(clk), .RN(rst), .Q(
        \regs[23][12] ) );
  DFFRHQX1 \regs_reg[23][11]  ( .D(n833), .CK(clk), .RN(rst), .Q(
        \regs[23][11] ) );
  DFFRHQX1 \regs_reg[23][10]  ( .D(n832), .CK(clk), .RN(rst), .Q(
        \regs[23][10] ) );
  DFFRHQX1 \regs_reg[23][9]  ( .D(n831), .CK(clk), .RN(rst), .Q(\regs[23][9] )
         );
  DFFRHQX1 \regs_reg[23][8]  ( .D(n830), .CK(clk), .RN(rst), .Q(\regs[23][8] )
         );
  DFFRHQX1 \regs_reg[23][7]  ( .D(n829), .CK(clk), .RN(rst), .Q(\regs[23][7] )
         );
  DFFRHQX1 \regs_reg[23][6]  ( .D(n828), .CK(clk), .RN(rst), .Q(\regs[23][6] )
         );
  DFFRHQX1 \regs_reg[23][5]  ( .D(n827), .CK(clk), .RN(rst), .Q(\regs[23][5] )
         );
  DFFRHQX1 \regs_reg[23][4]  ( .D(n826), .CK(clk), .RN(rst), .Q(\regs[23][4] )
         );
  DFFRHQX1 \regs_reg[23][3]  ( .D(n825), .CK(clk), .RN(rst), .Q(\regs[23][3] )
         );
  DFFRHQX1 \regs_reg[23][2]  ( .D(n824), .CK(clk), .RN(rst), .Q(\regs[23][2] )
         );
  DFFRHQX1 \regs_reg[23][1]  ( .D(n823), .CK(clk), .RN(rst), .Q(\regs[23][1] )
         );
  DFFRHQX1 \regs_reg[23][0]  ( .D(n822), .CK(clk), .RN(rst), .Q(\regs[23][0] )
         );
  DFFRHQX1 \regs_reg[19][31]  ( .D(n725), .CK(clk), .RN(rst), .Q(
        \regs[19][31] ) );
  DFFRHQX1 \regs_reg[19][30]  ( .D(n724), .CK(clk), .RN(rst), .Q(
        \regs[19][30] ) );
  DFFRHQX1 \regs_reg[19][29]  ( .D(n723), .CK(clk), .RN(rst), .Q(
        \regs[19][29] ) );
  DFFRHQX1 \regs_reg[19][28]  ( .D(n722), .CK(clk), .RN(rst), .Q(
        \regs[19][28] ) );
  DFFRHQX1 \regs_reg[19][27]  ( .D(n721), .CK(clk), .RN(rst), .Q(
        \regs[19][27] ) );
  DFFRHQX1 \regs_reg[19][26]  ( .D(n720), .CK(clk), .RN(rst), .Q(
        \regs[19][26] ) );
  DFFRHQX1 \regs_reg[19][25]  ( .D(n719), .CK(clk), .RN(rst), .Q(
        \regs[19][25] ) );
  DFFRHQX1 \regs_reg[19][24]  ( .D(n718), .CK(clk), .RN(rst), .Q(
        \regs[19][24] ) );
  DFFRHQX1 \regs_reg[19][15]  ( .D(n709), .CK(clk), .RN(rst), .Q(
        \regs[19][15] ) );
  DFFRHQX1 \regs_reg[19][14]  ( .D(n708), .CK(clk), .RN(rst), .Q(
        \regs[19][14] ) );
  DFFRHQX1 \regs_reg[19][13]  ( .D(n707), .CK(clk), .RN(rst), .Q(
        \regs[19][13] ) );
  DFFRHQX1 \regs_reg[19][12]  ( .D(n706), .CK(clk), .RN(rst), .Q(
        \regs[19][12] ) );
  DFFRHQX1 \regs_reg[19][11]  ( .D(n705), .CK(clk), .RN(rst), .Q(
        \regs[19][11] ) );
  DFFRHQX1 \regs_reg[19][10]  ( .D(n704), .CK(clk), .RN(rst), .Q(
        \regs[19][10] ) );
  DFFRHQX1 \regs_reg[19][9]  ( .D(n703), .CK(clk), .RN(rst), .Q(\regs[19][9] )
         );
  DFFRHQX1 \regs_reg[19][8]  ( .D(n702), .CK(clk), .RN(rst), .Q(\regs[19][8] )
         );
  DFFRHQX1 \regs_reg[19][7]  ( .D(n701), .CK(clk), .RN(rst), .Q(\regs[19][7] )
         );
  DFFRHQX1 \regs_reg[19][6]  ( .D(n700), .CK(clk), .RN(rst), .Q(\regs[19][6] )
         );
  DFFRHQX1 \regs_reg[19][5]  ( .D(n699), .CK(clk), .RN(rst), .Q(\regs[19][5] )
         );
  DFFRHQX1 \regs_reg[19][4]  ( .D(n698), .CK(clk), .RN(rst), .Q(\regs[19][4] )
         );
  DFFRHQX1 \regs_reg[19][3]  ( .D(n697), .CK(clk), .RN(rst), .Q(\regs[19][3] )
         );
  DFFRHQX1 \regs_reg[19][2]  ( .D(n696), .CK(clk), .RN(rst), .Q(\regs[19][2] )
         );
  DFFRHQX1 \regs_reg[19][1]  ( .D(n695), .CK(clk), .RN(rst), .Q(\regs[19][1] )
         );
  DFFRHQX1 \regs_reg[19][0]  ( .D(n694), .CK(clk), .RN(rst), .Q(\regs[19][0] )
         );
  DFFRHQX1 \regs_reg[15][31]  ( .D(n597), .CK(clk), .RN(rst), .Q(
        \regs[15][31] ) );
  DFFRHQX1 \regs_reg[15][30]  ( .D(n596), .CK(clk), .RN(rst), .Q(
        \regs[15][30] ) );
  DFFRHQX1 \regs_reg[15][29]  ( .D(n595), .CK(clk), .RN(rst), .Q(
        \regs[15][29] ) );
  DFFRHQX1 \regs_reg[15][28]  ( .D(n594), .CK(clk), .RN(rst), .Q(
        \regs[15][28] ) );
  DFFRHQX1 \regs_reg[15][27]  ( .D(n593), .CK(clk), .RN(rst), .Q(
        \regs[15][27] ) );
  DFFRHQX1 \regs_reg[15][26]  ( .D(n592), .CK(clk), .RN(rst), .Q(
        \regs[15][26] ) );
  DFFRHQX1 \regs_reg[15][25]  ( .D(n591), .CK(clk), .RN(rst), .Q(
        \regs[15][25] ) );
  DFFRHQX1 \regs_reg[15][24]  ( .D(n590), .CK(clk), .RN(rst), .Q(
        \regs[15][24] ) );
  DFFRHQX1 \regs_reg[15][15]  ( .D(n581), .CK(clk), .RN(rst), .Q(
        \regs[15][15] ) );
  DFFRHQX1 \regs_reg[15][14]  ( .D(n580), .CK(clk), .RN(rst), .Q(
        \regs[15][14] ) );
  DFFRHQX1 \regs_reg[15][13]  ( .D(n579), .CK(clk), .RN(rst), .Q(
        \regs[15][13] ) );
  DFFRHQX1 \regs_reg[15][12]  ( .D(n578), .CK(clk), .RN(rst), .Q(
        \regs[15][12] ) );
  DFFRHQX1 \regs_reg[15][11]  ( .D(n577), .CK(clk), .RN(rst), .Q(
        \regs[15][11] ) );
  DFFRHQX1 \regs_reg[15][10]  ( .D(n576), .CK(clk), .RN(rst), .Q(
        \regs[15][10] ) );
  DFFRHQX1 \regs_reg[15][9]  ( .D(n575), .CK(clk), .RN(rst), .Q(\regs[15][9] )
         );
  DFFRHQX1 \regs_reg[15][8]  ( .D(n574), .CK(clk), .RN(rst), .Q(\regs[15][8] )
         );
  DFFRHQX1 \regs_reg[15][7]  ( .D(n573), .CK(clk), .RN(rst), .Q(\regs[15][7] )
         );
  DFFRHQX1 \regs_reg[15][6]  ( .D(n572), .CK(clk), .RN(rst), .Q(\regs[15][6] )
         );
  DFFRHQX1 \regs_reg[15][5]  ( .D(n571), .CK(clk), .RN(rst), .Q(\regs[15][5] )
         );
  DFFRHQX1 \regs_reg[15][4]  ( .D(n570), .CK(clk), .RN(rst), .Q(\regs[15][4] )
         );
  DFFRHQX1 \regs_reg[15][3]  ( .D(n569), .CK(clk), .RN(rst), .Q(\regs[15][3] )
         );
  DFFRHQX1 \regs_reg[15][2]  ( .D(n568), .CK(clk), .RN(rst), .Q(\regs[15][2] )
         );
  DFFRHQX1 \regs_reg[15][1]  ( .D(n567), .CK(clk), .RN(rst), .Q(\regs[15][1] )
         );
  DFFRHQX1 \regs_reg[15][0]  ( .D(n566), .CK(clk), .RN(rst), .Q(\regs[15][0] )
         );
  DFFRHQX1 \regs_reg[11][31]  ( .D(n469), .CK(clk), .RN(rst), .Q(
        \regs[11][31] ) );
  DFFRHQX1 \regs_reg[11][30]  ( .D(n468), .CK(clk), .RN(rst), .Q(
        \regs[11][30] ) );
  DFFRHQX1 \regs_reg[11][29]  ( .D(n467), .CK(clk), .RN(rst), .Q(
        \regs[11][29] ) );
  DFFRHQX1 \regs_reg[11][28]  ( .D(n466), .CK(clk), .RN(rst), .Q(
        \regs[11][28] ) );
  DFFRHQX1 \regs_reg[11][27]  ( .D(n465), .CK(clk), .RN(rst), .Q(
        \regs[11][27] ) );
  DFFRHQX1 \regs_reg[11][26]  ( .D(n464), .CK(clk), .RN(rst), .Q(
        \regs[11][26] ) );
  DFFRHQX1 \regs_reg[11][25]  ( .D(n463), .CK(clk), .RN(rst), .Q(
        \regs[11][25] ) );
  DFFRHQX1 \regs_reg[11][24]  ( .D(n462), .CK(clk), .RN(rst), .Q(
        \regs[11][24] ) );
  DFFRHQX1 \regs_reg[11][15]  ( .D(n453), .CK(clk), .RN(rst), .Q(
        \regs[11][15] ) );
  DFFRHQX1 \regs_reg[11][14]  ( .D(n452), .CK(clk), .RN(rst), .Q(
        \regs[11][14] ) );
  DFFRHQX1 \regs_reg[11][13]  ( .D(n451), .CK(clk), .RN(rst), .Q(
        \regs[11][13] ) );
  DFFRHQX1 \regs_reg[11][12]  ( .D(n450), .CK(clk), .RN(rst), .Q(
        \regs[11][12] ) );
  DFFRHQX1 \regs_reg[11][11]  ( .D(n449), .CK(clk), .RN(rst), .Q(
        \regs[11][11] ) );
  DFFRHQX1 \regs_reg[11][10]  ( .D(n448), .CK(clk), .RN(rst), .Q(
        \regs[11][10] ) );
  DFFRHQX1 \regs_reg[11][9]  ( .D(n447), .CK(clk), .RN(rst), .Q(\regs[11][9] )
         );
  DFFRHQX1 \regs_reg[11][8]  ( .D(n446), .CK(clk), .RN(rst), .Q(\regs[11][8] )
         );
  DFFRHQX1 \regs_reg[11][7]  ( .D(n445), .CK(clk), .RN(rst), .Q(\regs[11][7] )
         );
  DFFRHQX1 \regs_reg[11][6]  ( .D(n444), .CK(clk), .RN(rst), .Q(\regs[11][6] )
         );
  DFFRHQX1 \regs_reg[11][5]  ( .D(n443), .CK(clk), .RN(rst), .Q(\regs[11][5] )
         );
  DFFRHQX1 \regs_reg[11][4]  ( .D(n442), .CK(clk), .RN(rst), .Q(\regs[11][4] )
         );
  DFFRHQX1 \regs_reg[11][3]  ( .D(n441), .CK(clk), .RN(rst), .Q(\regs[11][3] )
         );
  DFFRHQX1 \regs_reg[11][2]  ( .D(n440), .CK(clk), .RN(rst), .Q(\regs[11][2] )
         );
  DFFRHQX1 \regs_reg[11][1]  ( .D(n439), .CK(clk), .RN(rst), .Q(\regs[11][1] )
         );
  DFFRHQX1 \regs_reg[11][0]  ( .D(n438), .CK(clk), .RN(rst), .Q(\regs[11][0] )
         );
  DFFRHQX1 \regs_reg[7][31]  ( .D(n341), .CK(clk), .RN(rst), .Q(\regs[7][31] )
         );
  DFFRHQX1 \regs_reg[7][30]  ( .D(n340), .CK(clk), .RN(rst), .Q(\regs[7][30] )
         );
  DFFRHQX1 \regs_reg[7][29]  ( .D(n339), .CK(clk), .RN(rst), .Q(\regs[7][29] )
         );
  DFFRHQX1 \regs_reg[7][28]  ( .D(n338), .CK(clk), .RN(rst), .Q(\regs[7][28] )
         );
  DFFRHQX1 \regs_reg[7][27]  ( .D(n337), .CK(clk), .RN(rst), .Q(\regs[7][27] )
         );
  DFFRHQX1 \regs_reg[7][26]  ( .D(n336), .CK(clk), .RN(rst), .Q(\regs[7][26] )
         );
  DFFRHQX1 \regs_reg[7][25]  ( .D(n335), .CK(clk), .RN(rst), .Q(\regs[7][25] )
         );
  DFFRHQX1 \regs_reg[7][24]  ( .D(n334), .CK(clk), .RN(rst), .Q(\regs[7][24] )
         );
  DFFRHQX1 \regs_reg[7][15]  ( .D(n325), .CK(clk), .RN(rst), .Q(\regs[7][15] )
         );
  DFFRHQX1 \regs_reg[7][14]  ( .D(n324), .CK(clk), .RN(rst), .Q(\regs[7][14] )
         );
  DFFRHQX1 \regs_reg[7][13]  ( .D(n323), .CK(clk), .RN(rst), .Q(\regs[7][13] )
         );
  DFFRHQX1 \regs_reg[7][12]  ( .D(n322), .CK(clk), .RN(rst), .Q(\regs[7][12] )
         );
  DFFRHQX1 \regs_reg[7][11]  ( .D(n321), .CK(clk), .RN(rst), .Q(\regs[7][11] )
         );
  DFFRHQX1 \regs_reg[7][10]  ( .D(n320), .CK(clk), .RN(rst), .Q(\regs[7][10] )
         );
  DFFRHQX1 \regs_reg[7][9]  ( .D(n319), .CK(clk), .RN(rst), .Q(\regs[7][9] )
         );
  DFFRHQX1 \regs_reg[7][8]  ( .D(n318), .CK(clk), .RN(rst), .Q(\regs[7][8] )
         );
  DFFRHQX1 \regs_reg[7][7]  ( .D(n317), .CK(clk), .RN(rst), .Q(\regs[7][7] )
         );
  DFFRHQX1 \regs_reg[7][6]  ( .D(n316), .CK(clk), .RN(rst), .Q(\regs[7][6] )
         );
  DFFRHQX1 \regs_reg[7][5]  ( .D(n315), .CK(clk), .RN(rst), .Q(\regs[7][5] )
         );
  DFFRHQX1 \regs_reg[7][4]  ( .D(n314), .CK(clk), .RN(rst), .Q(\regs[7][4] )
         );
  DFFRHQX1 \regs_reg[7][3]  ( .D(n313), .CK(clk), .RN(rst), .Q(\regs[7][3] )
         );
  DFFRHQX1 \regs_reg[7][2]  ( .D(n312), .CK(clk), .RN(rst), .Q(\regs[7][2] )
         );
  DFFRHQX1 \regs_reg[7][1]  ( .D(n311), .CK(clk), .RN(rst), .Q(\regs[7][1] )
         );
  DFFRHQX1 \regs_reg[7][0]  ( .D(n310), .CK(clk), .RN(rst), .Q(\regs[7][0] )
         );
  DFFRHQX1 \regs_reg[3][31]  ( .D(n213), .CK(clk), .RN(rst), .Q(\regs[3][31] )
         );
  DFFRHQX1 \regs_reg[3][30]  ( .D(n212), .CK(clk), .RN(rst), .Q(\regs[3][30] )
         );
  DFFRHQX1 \regs_reg[3][29]  ( .D(n211), .CK(clk), .RN(rst), .Q(\regs[3][29] )
         );
  DFFRHQX1 \regs_reg[3][28]  ( .D(n210), .CK(clk), .RN(rst), .Q(\regs[3][28] )
         );
  DFFRHQX1 \regs_reg[3][27]  ( .D(n209), .CK(clk), .RN(rst), .Q(\regs[3][27] )
         );
  DFFRHQX1 \regs_reg[3][26]  ( .D(n208), .CK(clk), .RN(rst), .Q(\regs[3][26] )
         );
  DFFRHQX1 \regs_reg[3][25]  ( .D(n207), .CK(clk), .RN(rst), .Q(\regs[3][25] )
         );
  DFFRHQX1 \regs_reg[3][24]  ( .D(n206), .CK(clk), .RN(rst), .Q(\regs[3][24] )
         );
  DFFRHQX1 \regs_reg[3][19]  ( .D(n201), .CK(clk), .RN(rst), .Q(\regs[3][19] )
         );
  DFFRHQX1 \regs_reg[3][15]  ( .D(n197), .CK(clk), .RN(rst), .Q(\regs[3][15] )
         );
  DFFRHQX1 \regs_reg[3][14]  ( .D(n196), .CK(clk), .RN(rst), .Q(\regs[3][14] )
         );
  DFFRHQX1 \regs_reg[3][13]  ( .D(n195), .CK(clk), .RN(rst), .Q(\regs[3][13] )
         );
  DFFRHQX1 \regs_reg[3][12]  ( .D(n194), .CK(clk), .RN(rst), .Q(\regs[3][12] )
         );
  DFFRHQX1 \regs_reg[3][11]  ( .D(n193), .CK(clk), .RN(rst), .Q(\regs[3][11] )
         );
  DFFRHQX1 \regs_reg[3][10]  ( .D(n192), .CK(clk), .RN(rst), .Q(\regs[3][10] )
         );
  DFFRHQX1 \regs_reg[3][9]  ( .D(n191), .CK(clk), .RN(rst), .Q(\regs[3][9] )
         );
  DFFRHQX1 \regs_reg[3][8]  ( .D(n190), .CK(clk), .RN(rst), .Q(\regs[3][8] )
         );
  DFFRHQX1 \regs_reg[3][7]  ( .D(n189), .CK(clk), .RN(rst), .Q(\regs[3][7] )
         );
  DFFRHQX1 \regs_reg[3][6]  ( .D(n188), .CK(clk), .RN(rst), .Q(\regs[3][6] )
         );
  DFFRHQX1 \regs_reg[3][5]  ( .D(n187), .CK(clk), .RN(rst), .Q(\regs[3][5] )
         );
  DFFRHQX1 \regs_reg[3][4]  ( .D(n186), .CK(clk), .RN(rst), .Q(\regs[3][4] )
         );
  DFFRHQX1 \regs_reg[3][3]  ( .D(n185), .CK(clk), .RN(rst), .Q(\regs[3][3] )
         );
  DFFRHQX1 \regs_reg[3][2]  ( .D(n184), .CK(clk), .RN(rst), .Q(\regs[3][2] )
         );
  DFFRHQX1 \regs_reg[3][1]  ( .D(n183), .CK(clk), .RN(rst), .Q(\regs[3][1] )
         );
  DFFRHQX1 \regs_reg[3][0]  ( .D(n182), .CK(clk), .RN(rst), .Q(\regs[3][0] )
         );
  DFFRHQX1 \regs_reg[28][31]  ( .D(n1013), .CK(clk), .RN(rst), .Q(
        \regs[28][31] ) );
  DFFRHQX1 \regs_reg[28][30]  ( .D(n1012), .CK(clk), .RN(rst), .Q(
        \regs[28][30] ) );
  DFFRHQX1 \regs_reg[28][29]  ( .D(n1011), .CK(clk), .RN(rst), .Q(
        \regs[28][29] ) );
  DFFRHQX1 \regs_reg[28][28]  ( .D(n1010), .CK(clk), .RN(rst), .Q(
        \regs[28][28] ) );
  DFFRHQX1 \regs_reg[28][27]  ( .D(n1009), .CK(clk), .RN(rst), .Q(
        \regs[28][27] ) );
  DFFRHQX1 \regs_reg[28][26]  ( .D(n1008), .CK(clk), .RN(rst), .Q(
        \regs[28][26] ) );
  DFFRHQX1 \regs_reg[28][25]  ( .D(n1007), .CK(clk), .RN(rst), .Q(
        \regs[28][25] ) );
  DFFRHQX1 \regs_reg[28][24]  ( .D(n1006), .CK(clk), .RN(rst), .Q(
        \regs[28][24] ) );
  DFFRHQX1 \regs_reg[28][15]  ( .D(n997), .CK(clk), .RN(rst), .Q(
        \regs[28][15] ) );
  DFFRHQX1 \regs_reg[28][14]  ( .D(n996), .CK(clk), .RN(rst), .Q(
        \regs[28][14] ) );
  DFFRHQX1 \regs_reg[28][13]  ( .D(n995), .CK(clk), .RN(rst), .Q(
        \regs[28][13] ) );
  DFFRHQX1 \regs_reg[28][12]  ( .D(n994), .CK(clk), .RN(rst), .Q(
        \regs[28][12] ) );
  DFFRHQX1 \regs_reg[28][11]  ( .D(n993), .CK(clk), .RN(rst), .Q(
        \regs[28][11] ) );
  DFFRHQX1 \regs_reg[28][10]  ( .D(n992), .CK(clk), .RN(rst), .Q(
        \regs[28][10] ) );
  DFFRHQX1 \regs_reg[28][9]  ( .D(n991), .CK(clk), .RN(rst), .Q(\regs[28][9] )
         );
  DFFRHQX1 \regs_reg[28][8]  ( .D(n990), .CK(clk), .RN(rst), .Q(\regs[28][8] )
         );
  DFFRHQX1 \regs_reg[28][7]  ( .D(n989), .CK(clk), .RN(rst), .Q(\regs[28][7] )
         );
  DFFRHQX1 \regs_reg[28][6]  ( .D(n988), .CK(clk), .RN(rst), .Q(\regs[28][6] )
         );
  DFFRHQX1 \regs_reg[28][5]  ( .D(n987), .CK(clk), .RN(rst), .Q(\regs[28][5] )
         );
  DFFRHQX1 \regs_reg[28][4]  ( .D(n986), .CK(clk), .RN(rst), .Q(\regs[28][4] )
         );
  DFFRHQX1 \regs_reg[28][3]  ( .D(n985), .CK(clk), .RN(rst), .Q(\regs[28][3] )
         );
  DFFRHQX1 \regs_reg[28][2]  ( .D(n984), .CK(clk), .RN(rst), .Q(\regs[28][2] )
         );
  DFFRHQX1 \regs_reg[28][1]  ( .D(n983), .CK(clk), .RN(rst), .Q(\regs[28][1] )
         );
  DFFRHQX1 \regs_reg[28][0]  ( .D(n982), .CK(clk), .RN(rst), .Q(\regs[28][0] )
         );
  DFFRHQX1 \regs_reg[24][31]  ( .D(n885), .CK(clk), .RN(rst), .Q(
        \regs[24][31] ) );
  DFFRHQX1 \regs_reg[24][30]  ( .D(n884), .CK(clk), .RN(rst), .Q(
        \regs[24][30] ) );
  DFFRHQX1 \regs_reg[24][29]  ( .D(n883), .CK(clk), .RN(rst), .Q(
        \regs[24][29] ) );
  DFFRHQX1 \regs_reg[24][28]  ( .D(n882), .CK(clk), .RN(rst), .Q(
        \regs[24][28] ) );
  DFFRHQX1 \regs_reg[24][27]  ( .D(n881), .CK(clk), .RN(rst), .Q(
        \regs[24][27] ) );
  DFFRHQX1 \regs_reg[24][26]  ( .D(n880), .CK(clk), .RN(rst), .Q(
        \regs[24][26] ) );
  DFFRHQX1 \regs_reg[24][25]  ( .D(n879), .CK(clk), .RN(rst), .Q(
        \regs[24][25] ) );
  DFFRHQX1 \regs_reg[24][24]  ( .D(n878), .CK(clk), .RN(rst), .Q(
        \regs[24][24] ) );
  DFFRHQX1 \regs_reg[24][19]  ( .D(n873), .CK(clk), .RN(rst), .Q(
        \regs[24][19] ) );
  DFFRHQX1 \regs_reg[24][15]  ( .D(n869), .CK(clk), .RN(rst), .Q(
        \regs[24][15] ) );
  DFFRHQX1 \regs_reg[24][14]  ( .D(n868), .CK(clk), .RN(rst), .Q(
        \regs[24][14] ) );
  DFFRHQX1 \regs_reg[24][13]  ( .D(n867), .CK(clk), .RN(rst), .Q(
        \regs[24][13] ) );
  DFFRHQX1 \regs_reg[24][12]  ( .D(n866), .CK(clk), .RN(rst), .Q(
        \regs[24][12] ) );
  DFFRHQX1 \regs_reg[24][11]  ( .D(n865), .CK(clk), .RN(rst), .Q(
        \regs[24][11] ) );
  DFFRHQX1 \regs_reg[24][10]  ( .D(n864), .CK(clk), .RN(rst), .Q(
        \regs[24][10] ) );
  DFFRHQX1 \regs_reg[24][9]  ( .D(n863), .CK(clk), .RN(rst), .Q(\regs[24][9] )
         );
  DFFRHQX1 \regs_reg[24][8]  ( .D(n862), .CK(clk), .RN(rst), .Q(\regs[24][8] )
         );
  DFFRHQX1 \regs_reg[24][7]  ( .D(n861), .CK(clk), .RN(rst), .Q(\regs[24][7] )
         );
  DFFRHQX1 \regs_reg[24][6]  ( .D(n860), .CK(clk), .RN(rst), .Q(\regs[24][6] )
         );
  DFFRHQX1 \regs_reg[24][5]  ( .D(n859), .CK(clk), .RN(rst), .Q(\regs[24][5] )
         );
  DFFRHQX1 \regs_reg[24][4]  ( .D(n858), .CK(clk), .RN(rst), .Q(\regs[24][4] )
         );
  DFFRHQX1 \regs_reg[24][3]  ( .D(n857), .CK(clk), .RN(rst), .Q(\regs[24][3] )
         );
  DFFRHQX1 \regs_reg[24][2]  ( .D(n856), .CK(clk), .RN(rst), .Q(\regs[24][2] )
         );
  DFFRHQX1 \regs_reg[24][1]  ( .D(n855), .CK(clk), .RN(rst), .Q(\regs[24][1] )
         );
  DFFRHQX1 \regs_reg[24][0]  ( .D(n854), .CK(clk), .RN(rst), .Q(\regs[24][0] )
         );
  DFFRHQX1 \regs_reg[20][31]  ( .D(n757), .CK(clk), .RN(rst), .Q(
        \regs[20][31] ) );
  DFFRHQX1 \regs_reg[20][30]  ( .D(n756), .CK(clk), .RN(rst), .Q(
        \regs[20][30] ) );
  DFFRHQX1 \regs_reg[20][29]  ( .D(n755), .CK(clk), .RN(rst), .Q(
        \regs[20][29] ) );
  DFFRHQX1 \regs_reg[20][28]  ( .D(n754), .CK(clk), .RN(rst), .Q(
        \regs[20][28] ) );
  DFFRHQX1 \regs_reg[20][27]  ( .D(n753), .CK(clk), .RN(rst), .Q(
        \regs[20][27] ) );
  DFFRHQX1 \regs_reg[20][26]  ( .D(n752), .CK(clk), .RN(rst), .Q(
        \regs[20][26] ) );
  DFFRHQX1 \regs_reg[20][25]  ( .D(n751), .CK(clk), .RN(rst), .Q(
        \regs[20][25] ) );
  DFFRHQX1 \regs_reg[20][24]  ( .D(n750), .CK(clk), .RN(rst), .Q(
        \regs[20][24] ) );
  DFFRHQX1 \regs_reg[20][15]  ( .D(n741), .CK(clk), .RN(rst), .Q(
        \regs[20][15] ) );
  DFFRHQX1 \regs_reg[20][14]  ( .D(n740), .CK(clk), .RN(rst), .Q(
        \regs[20][14] ) );
  DFFRHQX1 \regs_reg[20][13]  ( .D(n739), .CK(clk), .RN(rst), .Q(
        \regs[20][13] ) );
  DFFRHQX1 \regs_reg[20][12]  ( .D(n738), .CK(clk), .RN(rst), .Q(
        \regs[20][12] ) );
  DFFRHQX1 \regs_reg[20][11]  ( .D(n737), .CK(clk), .RN(rst), .Q(
        \regs[20][11] ) );
  DFFRHQX1 \regs_reg[20][10]  ( .D(n736), .CK(clk), .RN(rst), .Q(
        \regs[20][10] ) );
  DFFRHQX1 \regs_reg[20][9]  ( .D(n735), .CK(clk), .RN(rst), .Q(\regs[20][9] )
         );
  DFFRHQX1 \regs_reg[20][8]  ( .D(n734), .CK(clk), .RN(rst), .Q(\regs[20][8] )
         );
  DFFRHQX1 \regs_reg[20][7]  ( .D(n733), .CK(clk), .RN(rst), .Q(\regs[20][7] )
         );
  DFFRHQX1 \regs_reg[20][6]  ( .D(n732), .CK(clk), .RN(rst), .Q(\regs[20][6] )
         );
  DFFRHQX1 \regs_reg[20][5]  ( .D(n731), .CK(clk), .RN(rst), .Q(\regs[20][5] )
         );
  DFFRHQX1 \regs_reg[20][4]  ( .D(n730), .CK(clk), .RN(rst), .Q(\regs[20][4] )
         );
  DFFRHQX1 \regs_reg[20][3]  ( .D(n729), .CK(clk), .RN(rst), .Q(\regs[20][3] )
         );
  DFFRHQX1 \regs_reg[20][2]  ( .D(n728), .CK(clk), .RN(rst), .Q(\regs[20][2] )
         );
  DFFRHQX1 \regs_reg[20][1]  ( .D(n727), .CK(clk), .RN(rst), .Q(\regs[20][1] )
         );
  DFFRHQX1 \regs_reg[20][0]  ( .D(n726), .CK(clk), .RN(rst), .Q(\regs[20][0] )
         );
  DFFRHQX1 \regs_reg[16][31]  ( .D(n629), .CK(clk), .RN(rst), .Q(
        \regs[16][31] ) );
  DFFRHQX1 \regs_reg[16][30]  ( .D(n628), .CK(clk), .RN(rst), .Q(
        \regs[16][30] ) );
  DFFRHQX1 \regs_reg[16][29]  ( .D(n627), .CK(clk), .RN(rst), .Q(
        \regs[16][29] ) );
  DFFRHQX1 \regs_reg[16][28]  ( .D(n626), .CK(clk), .RN(rst), .Q(
        \regs[16][28] ) );
  DFFRHQX1 \regs_reg[16][27]  ( .D(n625), .CK(clk), .RN(rst), .Q(
        \regs[16][27] ) );
  DFFRHQX1 \regs_reg[16][26]  ( .D(n624), .CK(clk), .RN(rst), .Q(
        \regs[16][26] ) );
  DFFRHQX1 \regs_reg[16][25]  ( .D(n623), .CK(clk), .RN(rst), .Q(
        \regs[16][25] ) );
  DFFRHQX1 \regs_reg[16][24]  ( .D(n622), .CK(clk), .RN(rst), .Q(
        \regs[16][24] ) );
  DFFRHQX1 \regs_reg[16][19]  ( .D(n617), .CK(clk), .RN(rst), .Q(
        \regs[16][19] ) );
  DFFRHQX1 \regs_reg[16][18]  ( .D(n616), .CK(clk), .RN(rst), .Q(
        \regs[16][18] ) );
  DFFRHQX1 \regs_reg[16][15]  ( .D(n613), .CK(clk), .RN(rst), .Q(
        \regs[16][15] ) );
  DFFRHQX1 \regs_reg[16][14]  ( .D(n612), .CK(clk), .RN(rst), .Q(
        \regs[16][14] ) );
  DFFRHQX1 \regs_reg[16][13]  ( .D(n611), .CK(clk), .RN(rst), .Q(
        \regs[16][13] ) );
  DFFRHQX1 \regs_reg[16][12]  ( .D(n610), .CK(clk), .RN(rst), .Q(
        \regs[16][12] ) );
  DFFRHQX1 \regs_reg[16][11]  ( .D(n609), .CK(clk), .RN(rst), .Q(
        \regs[16][11] ) );
  DFFRHQX1 \regs_reg[16][10]  ( .D(n608), .CK(clk), .RN(rst), .Q(
        \regs[16][10] ) );
  DFFRHQX1 \regs_reg[16][9]  ( .D(n607), .CK(clk), .RN(rst), .Q(\regs[16][9] )
         );
  DFFRHQX1 \regs_reg[16][8]  ( .D(n606), .CK(clk), .RN(rst), .Q(\regs[16][8] )
         );
  DFFRHQX1 \regs_reg[16][7]  ( .D(n605), .CK(clk), .RN(rst), .Q(\regs[16][7] )
         );
  DFFRHQX1 \regs_reg[16][6]  ( .D(n604), .CK(clk), .RN(rst), .Q(\regs[16][6] )
         );
  DFFRHQX1 \regs_reg[16][5]  ( .D(n603), .CK(clk), .RN(rst), .Q(\regs[16][5] )
         );
  DFFRHQX1 \regs_reg[16][4]  ( .D(n602), .CK(clk), .RN(rst), .Q(\regs[16][4] )
         );
  DFFRHQX1 \regs_reg[16][3]  ( .D(n601), .CK(clk), .RN(rst), .Q(\regs[16][3] )
         );
  DFFRHQX1 \regs_reg[16][2]  ( .D(n600), .CK(clk), .RN(rst), .Q(\regs[16][2] )
         );
  DFFRHQX1 \regs_reg[16][1]  ( .D(n599), .CK(clk), .RN(rst), .Q(\regs[16][1] )
         );
  DFFRHQX1 \regs_reg[16][0]  ( .D(n598), .CK(clk), .RN(rst), .Q(\regs[16][0] )
         );
  DFFRHQX1 \regs_reg[12][31]  ( .D(n501), .CK(clk), .RN(rst), .Q(
        \regs[12][31] ) );
  DFFRHQX1 \regs_reg[12][30]  ( .D(n500), .CK(clk), .RN(rst), .Q(
        \regs[12][30] ) );
  DFFRHQX1 \regs_reg[12][29]  ( .D(n499), .CK(clk), .RN(rst), .Q(
        \regs[12][29] ) );
  DFFRHQX1 \regs_reg[12][28]  ( .D(n498), .CK(clk), .RN(rst), .Q(
        \regs[12][28] ) );
  DFFRHQX1 \regs_reg[12][27]  ( .D(n497), .CK(clk), .RN(rst), .Q(
        \regs[12][27] ) );
  DFFRHQX1 \regs_reg[12][26]  ( .D(n496), .CK(clk), .RN(rst), .Q(
        \regs[12][26] ) );
  DFFRHQX1 \regs_reg[12][25]  ( .D(n495), .CK(clk), .RN(rst), .Q(
        \regs[12][25] ) );
  DFFRHQX1 \regs_reg[12][24]  ( .D(n494), .CK(clk), .RN(rst), .Q(
        \regs[12][24] ) );
  DFFRHQX1 \regs_reg[12][19]  ( .D(n489), .CK(clk), .RN(rst), .Q(
        \regs[12][19] ) );
  DFFRHQX1 \regs_reg[12][15]  ( .D(n485), .CK(clk), .RN(rst), .Q(
        \regs[12][15] ) );
  DFFRHQX1 \regs_reg[12][14]  ( .D(n484), .CK(clk), .RN(rst), .Q(
        \regs[12][14] ) );
  DFFRHQX1 \regs_reg[12][13]  ( .D(n483), .CK(clk), .RN(rst), .Q(
        \regs[12][13] ) );
  DFFRHQX1 \regs_reg[12][12]  ( .D(n482), .CK(clk), .RN(rst), .Q(
        \regs[12][12] ) );
  DFFRHQX1 \regs_reg[12][11]  ( .D(n481), .CK(clk), .RN(rst), .Q(
        \regs[12][11] ) );
  DFFRHQX1 \regs_reg[12][10]  ( .D(n480), .CK(clk), .RN(rst), .Q(
        \regs[12][10] ) );
  DFFRHQX1 \regs_reg[12][9]  ( .D(n479), .CK(clk), .RN(rst), .Q(\regs[12][9] )
         );
  DFFRHQX1 \regs_reg[12][8]  ( .D(n478), .CK(clk), .RN(rst), .Q(\regs[12][8] )
         );
  DFFRHQX1 \regs_reg[12][7]  ( .D(n477), .CK(clk), .RN(rst), .Q(\regs[12][7] )
         );
  DFFRHQX1 \regs_reg[12][6]  ( .D(n476), .CK(clk), .RN(rst), .Q(\regs[12][6] )
         );
  DFFRHQX1 \regs_reg[12][5]  ( .D(n475), .CK(clk), .RN(rst), .Q(\regs[12][5] )
         );
  DFFRHQX1 \regs_reg[12][4]  ( .D(n474), .CK(clk), .RN(rst), .Q(\regs[12][4] )
         );
  DFFRHQX1 \regs_reg[12][3]  ( .D(n473), .CK(clk), .RN(rst), .Q(\regs[12][3] )
         );
  DFFRHQX1 \regs_reg[12][2]  ( .D(n472), .CK(clk), .RN(rst), .Q(\regs[12][2] )
         );
  DFFRHQX1 \regs_reg[12][1]  ( .D(n471), .CK(clk), .RN(rst), .Q(\regs[12][1] )
         );
  DFFRHQX1 \regs_reg[12][0]  ( .D(n470), .CK(clk), .RN(rst), .Q(\regs[12][0] )
         );
  DFFRHQX1 \regs_reg[8][31]  ( .D(n373), .CK(clk), .RN(rst), .Q(\regs[8][31] )
         );
  DFFRHQX1 \regs_reg[8][30]  ( .D(n372), .CK(clk), .RN(rst), .Q(\regs[8][30] )
         );
  DFFRHQX1 \regs_reg[8][29]  ( .D(n371), .CK(clk), .RN(rst), .Q(\regs[8][29] )
         );
  DFFRHQX1 \regs_reg[8][28]  ( .D(n370), .CK(clk), .RN(rst), .Q(\regs[8][28] )
         );
  DFFRHQX1 \regs_reg[8][27]  ( .D(n369), .CK(clk), .RN(rst), .Q(\regs[8][27] )
         );
  DFFRHQX1 \regs_reg[8][26]  ( .D(n368), .CK(clk), .RN(rst), .Q(\regs[8][26] )
         );
  DFFRHQX1 \regs_reg[8][25]  ( .D(n367), .CK(clk), .RN(rst), .Q(\regs[8][25] )
         );
  DFFRHQX1 \regs_reg[8][24]  ( .D(n366), .CK(clk), .RN(rst), .Q(\regs[8][24] )
         );
  DFFRHQX1 \regs_reg[8][19]  ( .D(n361), .CK(clk), .RN(rst), .Q(\regs[8][19] )
         );
  DFFRHQX1 \regs_reg[8][18]  ( .D(n360), .CK(clk), .RN(rst), .Q(\regs[8][18] )
         );
  DFFRHQX1 \regs_reg[8][15]  ( .D(n357), .CK(clk), .RN(rst), .Q(\regs[8][15] )
         );
  DFFRHQX1 \regs_reg[8][14]  ( .D(n356), .CK(clk), .RN(rst), .Q(\regs[8][14] )
         );
  DFFRHQX1 \regs_reg[8][13]  ( .D(n355), .CK(clk), .RN(rst), .Q(\regs[8][13] )
         );
  DFFRHQX1 \regs_reg[8][12]  ( .D(n354), .CK(clk), .RN(rst), .Q(\regs[8][12] )
         );
  DFFRHQX1 \regs_reg[8][11]  ( .D(n353), .CK(clk), .RN(rst), .Q(\regs[8][11] )
         );
  DFFRHQX1 \regs_reg[8][10]  ( .D(n352), .CK(clk), .RN(rst), .Q(\regs[8][10] )
         );
  DFFRHQX1 \regs_reg[8][9]  ( .D(n351), .CK(clk), .RN(rst), .Q(\regs[8][9] )
         );
  DFFRHQX1 \regs_reg[8][8]  ( .D(n350), .CK(clk), .RN(rst), .Q(\regs[8][8] )
         );
  DFFRHQX1 \regs_reg[8][7]  ( .D(n349), .CK(clk), .RN(rst), .Q(\regs[8][7] )
         );
  DFFRHQX1 \regs_reg[8][6]  ( .D(n348), .CK(clk), .RN(rst), .Q(\regs[8][6] )
         );
  DFFRHQX1 \regs_reg[8][5]  ( .D(n347), .CK(clk), .RN(rst), .Q(\regs[8][5] )
         );
  DFFRHQX1 \regs_reg[8][4]  ( .D(n346), .CK(clk), .RN(rst), .Q(\regs[8][4] )
         );
  DFFRHQX1 \regs_reg[8][3]  ( .D(n345), .CK(clk), .RN(rst), .Q(\regs[8][3] )
         );
  DFFRHQX1 \regs_reg[8][2]  ( .D(n344), .CK(clk), .RN(rst), .Q(\regs[8][2] )
         );
  DFFRHQX1 \regs_reg[8][1]  ( .D(n343), .CK(clk), .RN(rst), .Q(\regs[8][1] )
         );
  DFFRHQX1 \regs_reg[8][0]  ( .D(n342), .CK(clk), .RN(rst), .Q(\regs[8][0] )
         );
  DFFRHQX1 \regs_reg[4][31]  ( .D(n245), .CK(clk), .RN(rst), .Q(\regs[4][31] )
         );
  DFFRHQX1 \regs_reg[4][30]  ( .D(n244), .CK(clk), .RN(rst), .Q(\regs[4][30] )
         );
  DFFRHQX1 \regs_reg[4][29]  ( .D(n243), .CK(clk), .RN(rst), .Q(\regs[4][29] )
         );
  DFFRHQX1 \regs_reg[4][28]  ( .D(n242), .CK(clk), .RN(rst), .Q(\regs[4][28] )
         );
  DFFRHQX1 \regs_reg[4][27]  ( .D(n241), .CK(clk), .RN(rst), .Q(\regs[4][27] )
         );
  DFFRHQX1 \regs_reg[4][26]  ( .D(n240), .CK(clk), .RN(rst), .Q(\regs[4][26] )
         );
  DFFRHQX1 \regs_reg[4][25]  ( .D(n239), .CK(clk), .RN(rst), .Q(\regs[4][25] )
         );
  DFFRHQX1 \regs_reg[4][24]  ( .D(n238), .CK(clk), .RN(rst), .Q(\regs[4][24] )
         );
  DFFRHQX1 \regs_reg[4][19]  ( .D(n233), .CK(clk), .RN(rst), .Q(\regs[4][19] )
         );
  DFFRHQX1 \regs_reg[4][18]  ( .D(n232), .CK(clk), .RN(rst), .Q(\regs[4][18] )
         );
  DFFRHQX1 \regs_reg[4][15]  ( .D(n229), .CK(clk), .RN(rst), .Q(\regs[4][15] )
         );
  DFFRHQX1 \regs_reg[4][14]  ( .D(n228), .CK(clk), .RN(rst), .Q(\regs[4][14] )
         );
  DFFRHQX1 \regs_reg[4][13]  ( .D(n227), .CK(clk), .RN(rst), .Q(\regs[4][13] )
         );
  DFFRHQX1 \regs_reg[4][12]  ( .D(n226), .CK(clk), .RN(rst), .Q(\regs[4][12] )
         );
  DFFRHQX1 \regs_reg[4][11]  ( .D(n225), .CK(clk), .RN(rst), .Q(\regs[4][11] )
         );
  DFFRHQX1 \regs_reg[4][10]  ( .D(n224), .CK(clk), .RN(rst), .Q(\regs[4][10] )
         );
  DFFRHQX1 \regs_reg[4][9]  ( .D(n223), .CK(clk), .RN(rst), .Q(\regs[4][9] )
         );
  DFFRHQX1 \regs_reg[4][8]  ( .D(n222), .CK(clk), .RN(rst), .Q(\regs[4][8] )
         );
  DFFRHQX1 \regs_reg[4][7]  ( .D(n221), .CK(clk), .RN(rst), .Q(\regs[4][7] )
         );
  DFFRHQX1 \regs_reg[4][6]  ( .D(n220), .CK(clk), .RN(rst), .Q(\regs[4][6] )
         );
  DFFRHQX1 \regs_reg[4][5]  ( .D(n219), .CK(clk), .RN(rst), .Q(\regs[4][5] )
         );
  DFFRHQX1 \regs_reg[4][4]  ( .D(n218), .CK(clk), .RN(rst), .Q(\regs[4][4] )
         );
  DFFRHQX1 \regs_reg[4][3]  ( .D(n217), .CK(clk), .RN(rst), .Q(\regs[4][3] )
         );
  DFFRHQX1 \regs_reg[4][2]  ( .D(n216), .CK(clk), .RN(rst), .Q(\regs[4][2] )
         );
  DFFRHQX1 \regs_reg[4][1]  ( .D(n215), .CK(clk), .RN(rst), .Q(\regs[4][1] )
         );
  DFFRHQX1 \regs_reg[4][0]  ( .D(n214), .CK(clk), .RN(rst), .Q(\regs[4][0] )
         );
  DFFRHQX1 \regs_reg[0][31]  ( .D(n117), .CK(clk), .RN(rst), .Q(\regs[0][31] )
         );
  DFFRHQX1 \regs_reg[0][30]  ( .D(n116), .CK(clk), .RN(rst), .Q(\regs[0][30] )
         );
  DFFRHQX1 \regs_reg[0][29]  ( .D(n115), .CK(clk), .RN(rst), .Q(\regs[0][29] )
         );
  DFFRHQX1 \regs_reg[0][28]  ( .D(n114), .CK(clk), .RN(rst), .Q(\regs[0][28] )
         );
  DFFRHQX1 \regs_reg[0][27]  ( .D(n113), .CK(clk), .RN(rst), .Q(\regs[0][27] )
         );
  DFFRHQX1 \regs_reg[0][26]  ( .D(n112), .CK(clk), .RN(rst), .Q(\regs[0][26] )
         );
  DFFRHQX1 \regs_reg[0][25]  ( .D(n111), .CK(clk), .RN(rst), .Q(\regs[0][25] )
         );
  DFFRHQX1 \regs_reg[0][24]  ( .D(n110), .CK(clk), .RN(rst), .Q(\regs[0][24] )
         );
  DFFRHQX1 \regs_reg[0][19]  ( .D(n105), .CK(clk), .RN(rst), .Q(\regs[0][19] )
         );
  DFFRHQX1 \regs_reg[0][18]  ( .D(n104), .CK(clk), .RN(rst), .Q(\regs[0][18] )
         );
  DFFRHQX1 \regs_reg[0][17]  ( .D(n103), .CK(clk), .RN(rst), .Q(\regs[0][17] )
         );
  DFFRHQX1 \regs_reg[0][16]  ( .D(n102), .CK(clk), .RN(rst), .Q(\regs[0][16] )
         );
  DFFRHQX1 \regs_reg[0][15]  ( .D(n101), .CK(clk), .RN(rst), .Q(\regs[0][15] )
         );
  DFFRHQX1 \regs_reg[0][14]  ( .D(n100), .CK(clk), .RN(rst), .Q(\regs[0][14] )
         );
  DFFRHQX1 \regs_reg[0][13]  ( .D(n99), .CK(clk), .RN(rst), .Q(\regs[0][13] )
         );
  DFFRHQX1 \regs_reg[0][12]  ( .D(n98), .CK(clk), .RN(rst), .Q(\regs[0][12] )
         );
  DFFRHQX1 \regs_reg[0][11]  ( .D(n97), .CK(clk), .RN(rst), .Q(\regs[0][11] )
         );
  DFFRHQX1 \regs_reg[0][10]  ( .D(n96), .CK(clk), .RN(rst), .Q(\regs[0][10] )
         );
  DFFRHQX1 \regs_reg[0][9]  ( .D(n95), .CK(clk), .RN(rst), .Q(\regs[0][9] ) );
  DFFRHQX1 \regs_reg[0][8]  ( .D(n94), .CK(clk), .RN(rst), .Q(\regs[0][8] ) );
  DFFRHQX1 \regs_reg[0][7]  ( .D(n93), .CK(clk), .RN(rst), .Q(\regs[0][7] ) );
  DFFRHQX1 \regs_reg[0][6]  ( .D(n92), .CK(clk), .RN(rst), .Q(\regs[0][6] ) );
  DFFRHQX1 \regs_reg[0][5]  ( .D(n91), .CK(clk), .RN(rst), .Q(\regs[0][5] ) );
  DFFRHQX1 \regs_reg[0][4]  ( .D(n90), .CK(clk), .RN(rst), .Q(\regs[0][4] ) );
  DFFRHQX1 \regs_reg[0][3]  ( .D(n89), .CK(clk), .RN(rst), .Q(\regs[0][3] ) );
  DFFRHQX1 \regs_reg[0][2]  ( .D(n88), .CK(clk), .RN(rst), .Q(\regs[0][2] ) );
  DFFRHQX1 \regs_reg[0][1]  ( .D(n87), .CK(clk), .RN(rst), .Q(\regs[0][1] ) );
  DFFRHQX1 \regs_reg[0][0]  ( .D(n86), .CK(clk), .RN(rst), .Q(\regs[0][0] ) );
  DFFRHQX1 \regs_reg[30][31]  ( .D(n1077), .CK(clk), .RN(rst), .Q(
        \regs[30][31] ) );
  DFFRHQX1 \regs_reg[30][30]  ( .D(n1076), .CK(clk), .RN(rst), .Q(
        \regs[30][30] ) );
  DFFRHQX1 \regs_reg[30][29]  ( .D(n1075), .CK(clk), .RN(rst), .Q(
        \regs[30][29] ) );
  DFFRHQX1 \regs_reg[30][28]  ( .D(n1074), .CK(clk), .RN(rst), .Q(
        \regs[30][28] ) );
  DFFRHQX1 \regs_reg[30][27]  ( .D(n1073), .CK(clk), .RN(rst), .Q(
        \regs[30][27] ) );
  DFFRHQX1 \regs_reg[30][26]  ( .D(n1072), .CK(clk), .RN(rst), .Q(
        \regs[30][26] ) );
  DFFRHQX1 \regs_reg[30][25]  ( .D(n1071), .CK(clk), .RN(rst), .Q(
        \regs[30][25] ) );
  DFFRHQX1 \regs_reg[30][24]  ( .D(n1070), .CK(clk), .RN(rst), .Q(
        \regs[30][24] ) );
  DFFRHQX1 \regs_reg[30][15]  ( .D(n1061), .CK(clk), .RN(rst), .Q(
        \regs[30][15] ) );
  DFFRHQX1 \regs_reg[30][14]  ( .D(n1060), .CK(clk), .RN(rst), .Q(
        \regs[30][14] ) );
  DFFRHQX1 \regs_reg[30][13]  ( .D(n1059), .CK(clk), .RN(rst), .Q(
        \regs[30][13] ) );
  DFFRHQX1 \regs_reg[30][12]  ( .D(n1058), .CK(clk), .RN(rst), .Q(
        \regs[30][12] ) );
  DFFRHQX1 \regs_reg[30][11]  ( .D(n1057), .CK(clk), .RN(rst), .Q(
        \regs[30][11] ) );
  DFFRHQX1 \regs_reg[30][10]  ( .D(n1056), .CK(clk), .RN(rst), .Q(
        \regs[30][10] ) );
  DFFRHQX1 \regs_reg[30][9]  ( .D(n1055), .CK(clk), .RN(rst), .Q(\regs[30][9] ) );
  DFFRHQX1 \regs_reg[30][8]  ( .D(n1054), .CK(clk), .RN(rst), .Q(\regs[30][8] ) );
  DFFRHQX1 \regs_reg[30][7]  ( .D(n1053), .CK(clk), .RN(rst), .Q(\regs[30][7] ) );
  DFFRHQX1 \regs_reg[30][6]  ( .D(n1052), .CK(clk), .RN(rst), .Q(\regs[30][6] ) );
  DFFRHQX1 \regs_reg[30][5]  ( .D(n1051), .CK(clk), .RN(rst), .Q(\regs[30][5] ) );
  DFFRHQX1 \regs_reg[30][4]  ( .D(n1050), .CK(clk), .RN(rst), .Q(\regs[30][4] ) );
  DFFRHQX1 \regs_reg[30][3]  ( .D(n1049), .CK(clk), .RN(rst), .Q(\regs[30][3] ) );
  DFFRHQX1 \regs_reg[30][2]  ( .D(n1048), .CK(clk), .RN(rst), .Q(\regs[30][2] ) );
  DFFRHQX1 \regs_reg[30][1]  ( .D(n1047), .CK(clk), .RN(rst), .Q(\regs[30][1] ) );
  DFFRHQX1 \regs_reg[30][0]  ( .D(n1046), .CK(clk), .RN(rst), .Q(\regs[30][0] ) );
  DFFRHQX1 \regs_reg[26][31]  ( .D(n949), .CK(clk), .RN(rst), .Q(
        \regs[26][31] ) );
  DFFRHQX1 \regs_reg[26][30]  ( .D(n948), .CK(clk), .RN(rst), .Q(
        \regs[26][30] ) );
  DFFRHQX1 \regs_reg[26][29]  ( .D(n947), .CK(clk), .RN(rst), .Q(
        \regs[26][29] ) );
  DFFRHQX1 \regs_reg[26][28]  ( .D(n946), .CK(clk), .RN(rst), .Q(
        \regs[26][28] ) );
  DFFRHQX1 \regs_reg[26][27]  ( .D(n945), .CK(clk), .RN(rst), .Q(
        \regs[26][27] ) );
  DFFRHQX1 \regs_reg[26][26]  ( .D(n944), .CK(clk), .RN(rst), .Q(
        \regs[26][26] ) );
  DFFRHQX1 \regs_reg[26][25]  ( .D(n943), .CK(clk), .RN(rst), .Q(
        \regs[26][25] ) );
  DFFRHQX1 \regs_reg[26][24]  ( .D(n942), .CK(clk), .RN(rst), .Q(
        \regs[26][24] ) );
  DFFRHQX1 \regs_reg[26][15]  ( .D(n933), .CK(clk), .RN(rst), .Q(
        \regs[26][15] ) );
  DFFRHQX1 \regs_reg[26][14]  ( .D(n932), .CK(clk), .RN(rst), .Q(
        \regs[26][14] ) );
  DFFRHQX1 \regs_reg[26][13]  ( .D(n931), .CK(clk), .RN(rst), .Q(
        \regs[26][13] ) );
  DFFRHQX1 \regs_reg[26][12]  ( .D(n930), .CK(clk), .RN(rst), .Q(
        \regs[26][12] ) );
  DFFRHQX1 \regs_reg[26][11]  ( .D(n929), .CK(clk), .RN(rst), .Q(
        \regs[26][11] ) );
  DFFRHQX1 \regs_reg[26][10]  ( .D(n928), .CK(clk), .RN(rst), .Q(
        \regs[26][10] ) );
  DFFRHQX1 \regs_reg[26][9]  ( .D(n927), .CK(clk), .RN(rst), .Q(\regs[26][9] )
         );
  DFFRHQX1 \regs_reg[26][8]  ( .D(n926), .CK(clk), .RN(rst), .Q(\regs[26][8] )
         );
  DFFRHQX1 \regs_reg[26][7]  ( .D(n925), .CK(clk), .RN(rst), .Q(\regs[26][7] )
         );
  DFFRHQX1 \regs_reg[26][6]  ( .D(n924), .CK(clk), .RN(rst), .Q(\regs[26][6] )
         );
  DFFRHQX1 \regs_reg[26][5]  ( .D(n923), .CK(clk), .RN(rst), .Q(\regs[26][5] )
         );
  DFFRHQX1 \regs_reg[26][4]  ( .D(n922), .CK(clk), .RN(rst), .Q(\regs[26][4] )
         );
  DFFRHQX1 \regs_reg[26][3]  ( .D(n921), .CK(clk), .RN(rst), .Q(\regs[26][3] )
         );
  DFFRHQX1 \regs_reg[26][2]  ( .D(n920), .CK(clk), .RN(rst), .Q(\regs[26][2] )
         );
  DFFRHQX1 \regs_reg[26][1]  ( .D(n919), .CK(clk), .RN(rst), .Q(\regs[26][1] )
         );
  DFFRHQX1 \regs_reg[26][0]  ( .D(n918), .CK(clk), .RN(rst), .Q(\regs[26][0] )
         );
  DFFRHQX1 \regs_reg[22][31]  ( .D(n821), .CK(clk), .RN(rst), .Q(
        \regs[22][31] ) );
  DFFRHQX1 \regs_reg[22][30]  ( .D(n820), .CK(clk), .RN(rst), .Q(
        \regs[22][30] ) );
  DFFRHQX1 \regs_reg[22][29]  ( .D(n819), .CK(clk), .RN(rst), .Q(
        \regs[22][29] ) );
  DFFRHQX1 \regs_reg[22][28]  ( .D(n818), .CK(clk), .RN(rst), .Q(
        \regs[22][28] ) );
  DFFRHQX1 \regs_reg[22][27]  ( .D(n817), .CK(clk), .RN(rst), .Q(
        \regs[22][27] ) );
  DFFRHQX1 \regs_reg[22][26]  ( .D(n816), .CK(clk), .RN(rst), .Q(
        \regs[22][26] ) );
  DFFRHQX1 \regs_reg[22][25]  ( .D(n815), .CK(clk), .RN(rst), .Q(
        \regs[22][25] ) );
  DFFRHQX1 \regs_reg[22][24]  ( .D(n814), .CK(clk), .RN(rst), .Q(
        \regs[22][24] ) );
  DFFRHQX1 \regs_reg[22][15]  ( .D(n805), .CK(clk), .RN(rst), .Q(
        \regs[22][15] ) );
  DFFRHQX1 \regs_reg[22][14]  ( .D(n804), .CK(clk), .RN(rst), .Q(
        \regs[22][14] ) );
  DFFRHQX1 \regs_reg[22][13]  ( .D(n803), .CK(clk), .RN(rst), .Q(
        \regs[22][13] ) );
  DFFRHQX1 \regs_reg[22][12]  ( .D(n802), .CK(clk), .RN(rst), .Q(
        \regs[22][12] ) );
  DFFRHQX1 \regs_reg[22][11]  ( .D(n801), .CK(clk), .RN(rst), .Q(
        \regs[22][11] ) );
  DFFRHQX1 \regs_reg[22][10]  ( .D(n800), .CK(clk), .RN(rst), .Q(
        \regs[22][10] ) );
  DFFRHQX1 \regs_reg[22][9]  ( .D(n799), .CK(clk), .RN(rst), .Q(\regs[22][9] )
         );
  DFFRHQX1 \regs_reg[22][8]  ( .D(n798), .CK(clk), .RN(rst), .Q(\regs[22][8] )
         );
  DFFRHQX1 \regs_reg[22][7]  ( .D(n797), .CK(clk), .RN(rst), .Q(\regs[22][7] )
         );
  DFFRHQX1 \regs_reg[22][6]  ( .D(n796), .CK(clk), .RN(rst), .Q(\regs[22][6] )
         );
  DFFRHQX1 \regs_reg[22][5]  ( .D(n795), .CK(clk), .RN(rst), .Q(\regs[22][5] )
         );
  DFFRHQX1 \regs_reg[22][4]  ( .D(n794), .CK(clk), .RN(rst), .Q(\regs[22][4] )
         );
  DFFRHQX1 \regs_reg[22][3]  ( .D(n793), .CK(clk), .RN(rst), .Q(\regs[22][3] )
         );
  DFFRHQX1 \regs_reg[22][2]  ( .D(n792), .CK(clk), .RN(rst), .Q(\regs[22][2] )
         );
  DFFRHQX1 \regs_reg[22][1]  ( .D(n791), .CK(clk), .RN(rst), .Q(\regs[22][1] )
         );
  DFFRHQX1 \regs_reg[22][0]  ( .D(n790), .CK(clk), .RN(rst), .Q(\regs[22][0] )
         );
  DFFRHQX1 \regs_reg[18][31]  ( .D(n693), .CK(clk), .RN(rst), .Q(
        \regs[18][31] ) );
  DFFRHQX1 \regs_reg[18][30]  ( .D(n692), .CK(clk), .RN(rst), .Q(
        \regs[18][30] ) );
  DFFRHQX1 \regs_reg[18][29]  ( .D(n691), .CK(clk), .RN(rst), .Q(
        \regs[18][29] ) );
  DFFRHQX1 \regs_reg[18][28]  ( .D(n690), .CK(clk), .RN(rst), .Q(
        \regs[18][28] ) );
  DFFRHQX1 \regs_reg[18][27]  ( .D(n689), .CK(clk), .RN(rst), .Q(
        \regs[18][27] ) );
  DFFRHQX1 \regs_reg[18][26]  ( .D(n688), .CK(clk), .RN(rst), .Q(
        \regs[18][26] ) );
  DFFRHQX1 \regs_reg[18][25]  ( .D(n687), .CK(clk), .RN(rst), .Q(
        \regs[18][25] ) );
  DFFRHQX1 \regs_reg[18][24]  ( .D(n686), .CK(clk), .RN(rst), .Q(
        \regs[18][24] ) );
  DFFRHQX1 \regs_reg[18][15]  ( .D(n677), .CK(clk), .RN(rst), .Q(
        \regs[18][15] ) );
  DFFRHQX1 \regs_reg[18][14]  ( .D(n676), .CK(clk), .RN(rst), .Q(
        \regs[18][14] ) );
  DFFRHQX1 \regs_reg[18][13]  ( .D(n675), .CK(clk), .RN(rst), .Q(
        \regs[18][13] ) );
  DFFRHQX1 \regs_reg[18][12]  ( .D(n674), .CK(clk), .RN(rst), .Q(
        \regs[18][12] ) );
  DFFRHQX1 \regs_reg[18][11]  ( .D(n673), .CK(clk), .RN(rst), .Q(
        \regs[18][11] ) );
  DFFRHQX1 \regs_reg[18][10]  ( .D(n672), .CK(clk), .RN(rst), .Q(
        \regs[18][10] ) );
  DFFRHQX1 \regs_reg[18][9]  ( .D(n671), .CK(clk), .RN(rst), .Q(\regs[18][9] )
         );
  DFFRHQX1 \regs_reg[18][8]  ( .D(n670), .CK(clk), .RN(rst), .Q(\regs[18][8] )
         );
  DFFRHQX1 \regs_reg[18][7]  ( .D(n669), .CK(clk), .RN(rst), .Q(\regs[18][7] )
         );
  DFFRHQX1 \regs_reg[18][6]  ( .D(n668), .CK(clk), .RN(rst), .Q(\regs[18][6] )
         );
  DFFRHQX1 \regs_reg[18][5]  ( .D(n667), .CK(clk), .RN(rst), .Q(\regs[18][5] )
         );
  DFFRHQX1 \regs_reg[18][4]  ( .D(n666), .CK(clk), .RN(rst), .Q(\regs[18][4] )
         );
  DFFRHQX1 \regs_reg[18][3]  ( .D(n665), .CK(clk), .RN(rst), .Q(\regs[18][3] )
         );
  DFFRHQX1 \regs_reg[18][2]  ( .D(n664), .CK(clk), .RN(rst), .Q(\regs[18][2] )
         );
  DFFRHQX1 \regs_reg[18][1]  ( .D(n663), .CK(clk), .RN(rst), .Q(\regs[18][1] )
         );
  DFFRHQX1 \regs_reg[18][0]  ( .D(n662), .CK(clk), .RN(rst), .Q(\regs[18][0] )
         );
  DFFRHQX1 \regs_reg[14][31]  ( .D(n565), .CK(clk), .RN(rst), .Q(
        \regs[14][31] ) );
  DFFRHQX1 \regs_reg[14][30]  ( .D(n564), .CK(clk), .RN(rst), .Q(
        \regs[14][30] ) );
  DFFRHQX1 \regs_reg[14][29]  ( .D(n563), .CK(clk), .RN(rst), .Q(
        \regs[14][29] ) );
  DFFRHQX1 \regs_reg[14][28]  ( .D(n562), .CK(clk), .RN(rst), .Q(
        \regs[14][28] ) );
  DFFRHQX1 \regs_reg[14][27]  ( .D(n561), .CK(clk), .RN(rst), .Q(
        \regs[14][27] ) );
  DFFRHQX1 \regs_reg[14][26]  ( .D(n560), .CK(clk), .RN(rst), .Q(
        \regs[14][26] ) );
  DFFRHQX1 \regs_reg[14][25]  ( .D(n559), .CK(clk), .RN(rst), .Q(
        \regs[14][25] ) );
  DFFRHQX1 \regs_reg[14][24]  ( .D(n558), .CK(clk), .RN(rst), .Q(
        \regs[14][24] ) );
  DFFRHQX1 \regs_reg[14][15]  ( .D(n549), .CK(clk), .RN(rst), .Q(
        \regs[14][15] ) );
  DFFRHQX1 \regs_reg[14][14]  ( .D(n548), .CK(clk), .RN(rst), .Q(
        \regs[14][14] ) );
  DFFRHQX1 \regs_reg[14][13]  ( .D(n547), .CK(clk), .RN(rst), .Q(
        \regs[14][13] ) );
  DFFRHQX1 \regs_reg[14][12]  ( .D(n546), .CK(clk), .RN(rst), .Q(
        \regs[14][12] ) );
  DFFRHQX1 \regs_reg[14][11]  ( .D(n545), .CK(clk), .RN(rst), .Q(
        \regs[14][11] ) );
  DFFRHQX1 \regs_reg[14][10]  ( .D(n544), .CK(clk), .RN(rst), .Q(
        \regs[14][10] ) );
  DFFRHQX1 \regs_reg[14][9]  ( .D(n543), .CK(clk), .RN(rst), .Q(\regs[14][9] )
         );
  DFFRHQX1 \regs_reg[14][8]  ( .D(n542), .CK(clk), .RN(rst), .Q(\regs[14][8] )
         );
  DFFRHQX1 \regs_reg[14][7]  ( .D(n541), .CK(clk), .RN(rst), .Q(\regs[14][7] )
         );
  DFFRHQX1 \regs_reg[14][6]  ( .D(n540), .CK(clk), .RN(rst), .Q(\regs[14][6] )
         );
  DFFRHQX1 \regs_reg[14][5]  ( .D(n539), .CK(clk), .RN(rst), .Q(\regs[14][5] )
         );
  DFFRHQX1 \regs_reg[14][4]  ( .D(n538), .CK(clk), .RN(rst), .Q(\regs[14][4] )
         );
  DFFRHQX1 \regs_reg[14][3]  ( .D(n537), .CK(clk), .RN(rst), .Q(\regs[14][3] )
         );
  DFFRHQX1 \regs_reg[14][2]  ( .D(n536), .CK(clk), .RN(rst), .Q(\regs[14][2] )
         );
  DFFRHQX1 \regs_reg[14][1]  ( .D(n535), .CK(clk), .RN(rst), .Q(\regs[14][1] )
         );
  DFFRHQX1 \regs_reg[14][0]  ( .D(n534), .CK(clk), .RN(rst), .Q(\regs[14][0] )
         );
  DFFRHQX1 \regs_reg[10][31]  ( .D(n437), .CK(clk), .RN(rst), .Q(
        \regs[10][31] ) );
  DFFRHQX1 \regs_reg[10][30]  ( .D(n436), .CK(clk), .RN(rst), .Q(
        \regs[10][30] ) );
  DFFRHQX1 \regs_reg[10][29]  ( .D(n435), .CK(clk), .RN(rst), .Q(
        \regs[10][29] ) );
  DFFRHQX1 \regs_reg[10][28]  ( .D(n434), .CK(clk), .RN(rst), .Q(
        \regs[10][28] ) );
  DFFRHQX1 \regs_reg[10][27]  ( .D(n433), .CK(clk), .RN(rst), .Q(
        \regs[10][27] ) );
  DFFRHQX1 \regs_reg[10][26]  ( .D(n432), .CK(clk), .RN(rst), .Q(
        \regs[10][26] ) );
  DFFRHQX1 \regs_reg[10][25]  ( .D(n431), .CK(clk), .RN(rst), .Q(
        \regs[10][25] ) );
  DFFRHQX1 \regs_reg[10][24]  ( .D(n430), .CK(clk), .RN(rst), .Q(
        \regs[10][24] ) );
  DFFRHQX1 \regs_reg[10][19]  ( .D(n425), .CK(clk), .RN(rst), .Q(
        \regs[10][19] ) );
  DFFRHQX1 \regs_reg[10][15]  ( .D(n421), .CK(clk), .RN(rst), .Q(
        \regs[10][15] ) );
  DFFRHQX1 \regs_reg[10][14]  ( .D(n420), .CK(clk), .RN(rst), .Q(
        \regs[10][14] ) );
  DFFRHQX1 \regs_reg[10][13]  ( .D(n419), .CK(clk), .RN(rst), .Q(
        \regs[10][13] ) );
  DFFRHQX1 \regs_reg[10][12]  ( .D(n418), .CK(clk), .RN(rst), .Q(
        \regs[10][12] ) );
  DFFRHQX1 \regs_reg[10][11]  ( .D(n417), .CK(clk), .RN(rst), .Q(
        \regs[10][11] ) );
  DFFRHQX1 \regs_reg[10][10]  ( .D(n416), .CK(clk), .RN(rst), .Q(
        \regs[10][10] ) );
  DFFRHQX1 \regs_reg[10][9]  ( .D(n415), .CK(clk), .RN(rst), .Q(\regs[10][9] )
         );
  DFFRHQX1 \regs_reg[10][8]  ( .D(n414), .CK(clk), .RN(rst), .Q(\regs[10][8] )
         );
  DFFRHQX1 \regs_reg[10][7]  ( .D(n413), .CK(clk), .RN(rst), .Q(\regs[10][7] )
         );
  DFFRHQX1 \regs_reg[10][6]  ( .D(n412), .CK(clk), .RN(rst), .Q(\regs[10][6] )
         );
  DFFRHQX1 \regs_reg[10][5]  ( .D(n411), .CK(clk), .RN(rst), .Q(\regs[10][5] )
         );
  DFFRHQX1 \regs_reg[10][4]  ( .D(n410), .CK(clk), .RN(rst), .Q(\regs[10][4] )
         );
  DFFRHQX1 \regs_reg[10][3]  ( .D(n409), .CK(clk), .RN(rst), .Q(\regs[10][3] )
         );
  DFFRHQX1 \regs_reg[10][2]  ( .D(n408), .CK(clk), .RN(rst), .Q(\regs[10][2] )
         );
  DFFRHQX1 \regs_reg[10][1]  ( .D(n407), .CK(clk), .RN(rst), .Q(\regs[10][1] )
         );
  DFFRHQX1 \regs_reg[10][0]  ( .D(n406), .CK(clk), .RN(rst), .Q(\regs[10][0] )
         );
  DFFRHQX1 \regs_reg[6][31]  ( .D(n309), .CK(clk), .RN(rst), .Q(\regs[6][31] )
         );
  DFFRHQX1 \regs_reg[6][30]  ( .D(n308), .CK(clk), .RN(rst), .Q(\regs[6][30] )
         );
  DFFRHQX1 \regs_reg[6][29]  ( .D(n307), .CK(clk), .RN(rst), .Q(\regs[6][29] )
         );
  DFFRHQX1 \regs_reg[6][28]  ( .D(n306), .CK(clk), .RN(rst), .Q(\regs[6][28] )
         );
  DFFRHQX1 \regs_reg[6][27]  ( .D(n305), .CK(clk), .RN(rst), .Q(\regs[6][27] )
         );
  DFFRHQX1 \regs_reg[6][26]  ( .D(n304), .CK(clk), .RN(rst), .Q(\regs[6][26] )
         );
  DFFRHQX1 \regs_reg[6][25]  ( .D(n303), .CK(clk), .RN(rst), .Q(\regs[6][25] )
         );
  DFFRHQX1 \regs_reg[6][24]  ( .D(n302), .CK(clk), .RN(rst), .Q(\regs[6][24] )
         );
  DFFRHQX1 \regs_reg[6][15]  ( .D(n293), .CK(clk), .RN(rst), .Q(\regs[6][15] )
         );
  DFFRHQX1 \regs_reg[6][14]  ( .D(n292), .CK(clk), .RN(rst), .Q(\regs[6][14] )
         );
  DFFRHQX1 \regs_reg[6][13]  ( .D(n291), .CK(clk), .RN(rst), .Q(\regs[6][13] )
         );
  DFFRHQX1 \regs_reg[6][12]  ( .D(n290), .CK(clk), .RN(rst), .Q(\regs[6][12] )
         );
  DFFRHQX1 \regs_reg[6][11]  ( .D(n289), .CK(clk), .RN(rst), .Q(\regs[6][11] )
         );
  DFFRHQX1 \regs_reg[6][10]  ( .D(n288), .CK(clk), .RN(rst), .Q(\regs[6][10] )
         );
  DFFRHQX1 \regs_reg[6][9]  ( .D(n287), .CK(clk), .RN(rst), .Q(\regs[6][9] )
         );
  DFFRHQX1 \regs_reg[6][8]  ( .D(n286), .CK(clk), .RN(rst), .Q(\regs[6][8] )
         );
  DFFRHQX1 \regs_reg[6][7]  ( .D(n285), .CK(clk), .RN(rst), .Q(\regs[6][7] )
         );
  DFFRHQX1 \regs_reg[6][6]  ( .D(n284), .CK(clk), .RN(rst), .Q(\regs[6][6] )
         );
  DFFRHQX1 \regs_reg[6][5]  ( .D(n283), .CK(clk), .RN(rst), .Q(\regs[6][5] )
         );
  DFFRHQX1 \regs_reg[6][4]  ( .D(n282), .CK(clk), .RN(rst), .Q(\regs[6][4] )
         );
  DFFRHQX1 \regs_reg[6][3]  ( .D(n281), .CK(clk), .RN(rst), .Q(\regs[6][3] )
         );
  DFFRHQX1 \regs_reg[6][2]  ( .D(n280), .CK(clk), .RN(rst), .Q(\regs[6][2] )
         );
  DFFRHQX1 \regs_reg[6][1]  ( .D(n279), .CK(clk), .RN(rst), .Q(\regs[6][1] )
         );
  DFFRHQX1 \regs_reg[6][0]  ( .D(n278), .CK(clk), .RN(rst), .Q(\regs[6][0] )
         );
  DFFRHQX1 \regs_reg[2][31]  ( .D(n181), .CK(clk), .RN(rst), .Q(\regs[2][31] )
         );
  DFFRHQX1 \regs_reg[2][30]  ( .D(n180), .CK(clk), .RN(rst), .Q(\regs[2][30] )
         );
  DFFRHQX1 \regs_reg[2][29]  ( .D(n179), .CK(clk), .RN(rst), .Q(\regs[2][29] )
         );
  DFFRHQX1 \regs_reg[2][28]  ( .D(n178), .CK(clk), .RN(rst), .Q(\regs[2][28] )
         );
  DFFRHQX1 \regs_reg[2][27]  ( .D(n177), .CK(clk), .RN(rst), .Q(\regs[2][27] )
         );
  DFFRHQX1 \regs_reg[2][26]  ( .D(n176), .CK(clk), .RN(rst), .Q(\regs[2][26] )
         );
  DFFRHQX1 \regs_reg[2][25]  ( .D(n175), .CK(clk), .RN(rst), .Q(\regs[2][25] )
         );
  DFFRHQX1 \regs_reg[2][24]  ( .D(n174), .CK(clk), .RN(rst), .Q(\regs[2][24] )
         );
  DFFRHQX1 \regs_reg[2][19]  ( .D(n169), .CK(clk), .RN(rst), .Q(\regs[2][19] )
         );
  DFFRHQX1 \regs_reg[2][18]  ( .D(n168), .CK(clk), .RN(rst), .Q(\regs[2][18] )
         );
  DFFRHQX1 \regs_reg[2][15]  ( .D(n165), .CK(clk), .RN(rst), .Q(\regs[2][15] )
         );
  DFFRHQX1 \regs_reg[2][14]  ( .D(n164), .CK(clk), .RN(rst), .Q(\regs[2][14] )
         );
  DFFRHQX1 \regs_reg[2][13]  ( .D(n163), .CK(clk), .RN(rst), .Q(\regs[2][13] )
         );
  DFFRHQX1 \regs_reg[2][12]  ( .D(n162), .CK(clk), .RN(rst), .Q(\regs[2][12] )
         );
  DFFRHQX1 \regs_reg[2][11]  ( .D(n161), .CK(clk), .RN(rst), .Q(\regs[2][11] )
         );
  DFFRHQX1 \regs_reg[2][10]  ( .D(n160), .CK(clk), .RN(rst), .Q(\regs[2][10] )
         );
  DFFRHQX1 \regs_reg[2][9]  ( .D(n159), .CK(clk), .RN(rst), .Q(\regs[2][9] )
         );
  DFFRHQX1 \regs_reg[2][8]  ( .D(n158), .CK(clk), .RN(rst), .Q(\regs[2][8] )
         );
  DFFRHQX1 \regs_reg[2][7]  ( .D(n157), .CK(clk), .RN(rst), .Q(\regs[2][7] )
         );
  DFFRHQX1 \regs_reg[2][6]  ( .D(n156), .CK(clk), .RN(rst), .Q(\regs[2][6] )
         );
  DFFRHQX1 \regs_reg[2][5]  ( .D(n155), .CK(clk), .RN(rst), .Q(\regs[2][5] )
         );
  DFFRHQX1 \regs_reg[2][4]  ( .D(n154), .CK(clk), .RN(rst), .Q(\regs[2][4] )
         );
  DFFRHQX1 \regs_reg[2][3]  ( .D(n153), .CK(clk), .RN(rst), .Q(\regs[2][3] )
         );
  DFFRHQX1 \regs_reg[2][2]  ( .D(n152), .CK(clk), .RN(rst), .Q(\regs[2][2] )
         );
  DFFRHQX1 \regs_reg[2][1]  ( .D(n151), .CK(clk), .RN(rst), .Q(\regs[2][1] )
         );
  DFFRHQX1 \regs_reg[2][0]  ( .D(n150), .CK(clk), .RN(rst), .Q(\regs[2][0] )
         );
  DFFRHQX1 \regs_reg[29][23]  ( .D(n1037), .CK(clk), .RN(rst), .Q(
        \regs[29][23] ) );
  DFFRHQX1 \regs_reg[29][22]  ( .D(n1036), .CK(clk), .RN(rst), .Q(
        \regs[29][22] ) );
  DFFRHQX1 \regs_reg[29][21]  ( .D(n1035), .CK(clk), .RN(rst), .Q(
        \regs[29][21] ) );
  DFFRHQX1 \regs_reg[29][20]  ( .D(n1034), .CK(clk), .RN(rst), .Q(
        \regs[29][20] ) );
  DFFRHQX1 \regs_reg[29][19]  ( .D(n1033), .CK(clk), .RN(rst), .Q(
        \regs[29][19] ) );
  DFFRHQX1 \regs_reg[29][18]  ( .D(n1032), .CK(clk), .RN(rst), .Q(
        \regs[29][18] ) );
  DFFRHQX1 \regs_reg[29][17]  ( .D(n1031), .CK(clk), .RN(rst), .Q(
        \regs[29][17] ) );
  DFFRHQX1 \regs_reg[29][16]  ( .D(n1030), .CK(clk), .RN(rst), .Q(
        \regs[29][16] ) );
  DFFRHQX1 \regs_reg[25][23]  ( .D(n909), .CK(clk), .RN(rst), .Q(
        \regs[25][23] ) );
  DFFRHQX1 \regs_reg[25][22]  ( .D(n908), .CK(clk), .RN(rst), .Q(
        \regs[25][22] ) );
  DFFRHQX1 \regs_reg[25][21]  ( .D(n907), .CK(clk), .RN(rst), .Q(
        \regs[25][21] ) );
  DFFRHQX1 \regs_reg[25][20]  ( .D(n906), .CK(clk), .RN(rst), .Q(
        \regs[25][20] ) );
  DFFRHQX1 \regs_reg[25][19]  ( .D(n905), .CK(clk), .RN(rst), .Q(
        \regs[25][19] ) );
  DFFRHQX1 \regs_reg[25][18]  ( .D(n904), .CK(clk), .RN(rst), .Q(
        \regs[25][18] ) );
  DFFRHQX1 \regs_reg[25][17]  ( .D(n903), .CK(clk), .RN(rst), .Q(
        \regs[25][17] ) );
  DFFRHQX1 \regs_reg[25][16]  ( .D(n902), .CK(clk), .RN(rst), .Q(
        \regs[25][16] ) );
  DFFRHQX1 \regs_reg[21][23]  ( .D(n781), .CK(clk), .RN(rst), .Q(
        \regs[21][23] ) );
  DFFRHQX1 \regs_reg[21][22]  ( .D(n780), .CK(clk), .RN(rst), .Q(
        \regs[21][22] ) );
  DFFRHQX1 \regs_reg[21][21]  ( .D(n779), .CK(clk), .RN(rst), .Q(
        \regs[21][21] ) );
  DFFRHQX1 \regs_reg[21][20]  ( .D(n778), .CK(clk), .RN(rst), .Q(
        \regs[21][20] ) );
  DFFRHQX1 \regs_reg[21][19]  ( .D(n777), .CK(clk), .RN(rst), .Q(
        \regs[21][19] ) );
  DFFRHQX1 \regs_reg[21][18]  ( .D(n776), .CK(clk), .RN(rst), .Q(
        \regs[21][18] ) );
  DFFRHQX1 \regs_reg[21][17]  ( .D(n775), .CK(clk), .RN(rst), .Q(
        \regs[21][17] ) );
  DFFRHQX1 \regs_reg[21][16]  ( .D(n774), .CK(clk), .RN(rst), .Q(
        \regs[21][16] ) );
  DFFRHQX1 \regs_reg[17][23]  ( .D(n653), .CK(clk), .RN(rst), .Q(
        \regs[17][23] ) );
  DFFRHQX1 \regs_reg[17][22]  ( .D(n652), .CK(clk), .RN(rst), .Q(
        \regs[17][22] ) );
  DFFRHQX1 \regs_reg[17][21]  ( .D(n651), .CK(clk), .RN(rst), .Q(
        \regs[17][21] ) );
  DFFRHQX1 \regs_reg[17][20]  ( .D(n650), .CK(clk), .RN(rst), .Q(
        \regs[17][20] ) );
  DFFRHQX1 \regs_reg[17][18]  ( .D(n648), .CK(clk), .RN(rst), .Q(
        \regs[17][18] ) );
  DFFRHQX1 \regs_reg[17][17]  ( .D(n647), .CK(clk), .RN(rst), .Q(
        \regs[17][17] ) );
  DFFRHQX1 \regs_reg[17][16]  ( .D(n646), .CK(clk), .RN(rst), .Q(
        \regs[17][16] ) );
  DFFRHQX1 \regs_reg[13][23]  ( .D(n525), .CK(clk), .RN(rst), .Q(
        \regs[13][23] ) );
  DFFRHQX1 \regs_reg[13][22]  ( .D(n524), .CK(clk), .RN(rst), .Q(
        \regs[13][22] ) );
  DFFRHQX1 \regs_reg[13][21]  ( .D(n523), .CK(clk), .RN(rst), .Q(
        \regs[13][21] ) );
  DFFRHQX1 \regs_reg[13][20]  ( .D(n522), .CK(clk), .RN(rst), .Q(
        \regs[13][20] ) );
  DFFRHQX1 \regs_reg[13][19]  ( .D(n521), .CK(clk), .RN(rst), .Q(
        \regs[13][19] ) );
  DFFRHQX1 \regs_reg[13][18]  ( .D(n520), .CK(clk), .RN(rst), .Q(
        \regs[13][18] ) );
  DFFRHQX1 \regs_reg[13][17]  ( .D(n519), .CK(clk), .RN(rst), .Q(
        \regs[13][17] ) );
  DFFRHQX1 \regs_reg[13][16]  ( .D(n518), .CK(clk), .RN(rst), .Q(
        \regs[13][16] ) );
  DFFRHQX1 \regs_reg[9][23]  ( .D(n397), .CK(clk), .RN(rst), .Q(\regs[9][23] )
         );
  DFFRHQX1 \regs_reg[9][22]  ( .D(n396), .CK(clk), .RN(rst), .Q(\regs[9][22] )
         );
  DFFRHQX1 \regs_reg[9][21]  ( .D(n395), .CK(clk), .RN(rst), .Q(\regs[9][21] )
         );
  DFFRHQX1 \regs_reg[9][20]  ( .D(n394), .CK(clk), .RN(rst), .Q(\regs[9][20] )
         );
  DFFRHQX1 \regs_reg[9][18]  ( .D(n392), .CK(clk), .RN(rst), .Q(\regs[9][18] )
         );
  DFFRHQX1 \regs_reg[9][17]  ( .D(n391), .CK(clk), .RN(rst), .Q(\regs[9][17] )
         );
  DFFRHQX1 \regs_reg[9][16]  ( .D(n390), .CK(clk), .RN(rst), .Q(\regs[9][16] )
         );
  DFFRHQX1 \regs_reg[5][23]  ( .D(n269), .CK(clk), .RN(rst), .Q(\regs[5][23] )
         );
  DFFRHQX1 \regs_reg[5][22]  ( .D(n268), .CK(clk), .RN(rst), .Q(\regs[5][22] )
         );
  DFFRHQX1 \regs_reg[5][21]  ( .D(n267), .CK(clk), .RN(rst), .Q(\regs[5][21] )
         );
  DFFRHQX1 \regs_reg[5][20]  ( .D(n266), .CK(clk), .RN(rst), .Q(\regs[5][20] )
         );
  DFFRHQX1 \regs_reg[5][18]  ( .D(n264), .CK(clk), .RN(rst), .Q(\regs[5][18] )
         );
  DFFRHQX1 \regs_reg[5][17]  ( .D(n263), .CK(clk), .RN(rst), .Q(\regs[5][17] )
         );
  DFFRHQX1 \regs_reg[5][16]  ( .D(n262), .CK(clk), .RN(rst), .Q(\regs[5][16] )
         );
  DFFRHQX1 \regs_reg[1][23]  ( .D(n141), .CK(clk), .RN(rst), .Q(\regs[1][23] )
         );
  DFFRHQX1 \regs_reg[1][22]  ( .D(n140), .CK(clk), .RN(rst), .Q(\regs[1][22] )
         );
  DFFRHQX1 \regs_reg[1][21]  ( .D(n139), .CK(clk), .RN(rst), .Q(\regs[1][21] )
         );
  DFFRHQX1 \regs_reg[1][20]  ( .D(n138), .CK(clk), .RN(rst), .Q(\regs[1][20] )
         );
  DFFRHQX1 \regs_reg[1][17]  ( .D(n135), .CK(clk), .RN(rst), .Q(\regs[1][17] )
         );
  DFFRHQX1 \regs_reg[1][16]  ( .D(n134), .CK(clk), .RN(rst), .Q(\regs[1][16] )
         );
  DFFRHQX1 \regs_reg[31][23]  ( .D(n1101), .CK(clk), .RN(rst), .Q(
        \regs[31][23] ) );
  DFFRHQX1 \regs_reg[31][22]  ( .D(n1100), .CK(clk), .RN(rst), .Q(
        \regs[31][22] ) );
  DFFRHQX1 \regs_reg[31][21]  ( .D(n1099), .CK(clk), .RN(rst), .Q(
        \regs[31][21] ) );
  DFFRHQX1 \regs_reg[31][20]  ( .D(n1098), .CK(clk), .RN(rst), .Q(
        \regs[31][20] ) );
  DFFRHQX1 \regs_reg[31][19]  ( .D(n1097), .CK(clk), .RN(rst), .Q(
        \regs[31][19] ) );
  DFFRHQX1 \regs_reg[31][18]  ( .D(n1096), .CK(clk), .RN(rst), .Q(
        \regs[31][18] ) );
  DFFRHQX1 \regs_reg[31][17]  ( .D(n1095), .CK(clk), .RN(rst), .Q(
        \regs[31][17] ) );
  DFFRHQX1 \regs_reg[31][16]  ( .D(n1094), .CK(clk), .RN(rst), .Q(
        \regs[31][16] ) );
  DFFRHQX1 \regs_reg[27][23]  ( .D(n973), .CK(clk), .RN(rst), .Q(
        \regs[27][23] ) );
  DFFRHQX1 \regs_reg[27][22]  ( .D(n972), .CK(clk), .RN(rst), .Q(
        \regs[27][22] ) );
  DFFRHQX1 \regs_reg[27][21]  ( .D(n971), .CK(clk), .RN(rst), .Q(
        \regs[27][21] ) );
  DFFRHQX1 \regs_reg[27][20]  ( .D(n970), .CK(clk), .RN(rst), .Q(
        \regs[27][20] ) );
  DFFRHQX1 \regs_reg[27][19]  ( .D(n969), .CK(clk), .RN(rst), .Q(
        \regs[27][19] ) );
  DFFRHQX1 \regs_reg[27][18]  ( .D(n968), .CK(clk), .RN(rst), .Q(
        \regs[27][18] ) );
  DFFRHQX1 \regs_reg[27][17]  ( .D(n967), .CK(clk), .RN(rst), .Q(
        \regs[27][17] ) );
  DFFRHQX1 \regs_reg[27][16]  ( .D(n966), .CK(clk), .RN(rst), .Q(
        \regs[27][16] ) );
  DFFRHQX1 \regs_reg[23][23]  ( .D(n845), .CK(clk), .RN(rst), .Q(
        \regs[23][23] ) );
  DFFRHQX1 \regs_reg[23][22]  ( .D(n844), .CK(clk), .RN(rst), .Q(
        \regs[23][22] ) );
  DFFRHQX1 \regs_reg[23][21]  ( .D(n843), .CK(clk), .RN(rst), .Q(
        \regs[23][21] ) );
  DFFRHQX1 \regs_reg[23][20]  ( .D(n842), .CK(clk), .RN(rst), .Q(
        \regs[23][20] ) );
  DFFRHQX1 \regs_reg[23][19]  ( .D(n841), .CK(clk), .RN(rst), .Q(
        \regs[23][19] ) );
  DFFRHQX1 \regs_reg[23][18]  ( .D(n840), .CK(clk), .RN(rst), .Q(
        \regs[23][18] ) );
  DFFRHQX1 \regs_reg[23][17]  ( .D(n839), .CK(clk), .RN(rst), .Q(
        \regs[23][17] ) );
  DFFRHQX1 \regs_reg[23][16]  ( .D(n838), .CK(clk), .RN(rst), .Q(
        \regs[23][16] ) );
  DFFRHQX1 \regs_reg[19][23]  ( .D(n717), .CK(clk), .RN(rst), .Q(
        \regs[19][23] ) );
  DFFRHQX1 \regs_reg[19][22]  ( .D(n716), .CK(clk), .RN(rst), .Q(
        \regs[19][22] ) );
  DFFRHQX1 \regs_reg[19][21]  ( .D(n715), .CK(clk), .RN(rst), .Q(
        \regs[19][21] ) );
  DFFRHQX1 \regs_reg[19][20]  ( .D(n714), .CK(clk), .RN(rst), .Q(
        \regs[19][20] ) );
  DFFRHQX1 \regs_reg[19][19]  ( .D(n713), .CK(clk), .RN(rst), .Q(
        \regs[19][19] ) );
  DFFRHQX1 \regs_reg[19][18]  ( .D(n712), .CK(clk), .RN(rst), .Q(
        \regs[19][18] ) );
  DFFRHQX1 \regs_reg[19][17]  ( .D(n711), .CK(clk), .RN(rst), .Q(
        \regs[19][17] ) );
  DFFRHQX1 \regs_reg[19][16]  ( .D(n710), .CK(clk), .RN(rst), .Q(
        \regs[19][16] ) );
  DFFRHQX1 \regs_reg[15][23]  ( .D(n589), .CK(clk), .RN(rst), .Q(
        \regs[15][23] ) );
  DFFRHQX1 \regs_reg[15][22]  ( .D(n588), .CK(clk), .RN(rst), .Q(
        \regs[15][22] ) );
  DFFRHQX1 \regs_reg[15][21]  ( .D(n587), .CK(clk), .RN(rst), .Q(
        \regs[15][21] ) );
  DFFRHQX1 \regs_reg[15][20]  ( .D(n586), .CK(clk), .RN(rst), .Q(
        \regs[15][20] ) );
  DFFRHQX1 \regs_reg[15][19]  ( .D(n585), .CK(clk), .RN(rst), .Q(
        \regs[15][19] ) );
  DFFRHQX1 \regs_reg[15][18]  ( .D(n584), .CK(clk), .RN(rst), .Q(
        \regs[15][18] ) );
  DFFRHQX1 \regs_reg[15][17]  ( .D(n583), .CK(clk), .RN(rst), .Q(
        \regs[15][17] ) );
  DFFRHQX1 \regs_reg[15][16]  ( .D(n582), .CK(clk), .RN(rst), .Q(
        \regs[15][16] ) );
  DFFRHQX1 \regs_reg[11][23]  ( .D(n461), .CK(clk), .RN(rst), .Q(
        \regs[11][23] ) );
  DFFRHQX1 \regs_reg[11][22]  ( .D(n460), .CK(clk), .RN(rst), .Q(
        \regs[11][22] ) );
  DFFRHQX1 \regs_reg[11][21]  ( .D(n459), .CK(clk), .RN(rst), .Q(
        \regs[11][21] ) );
  DFFRHQX1 \regs_reg[11][20]  ( .D(n458), .CK(clk), .RN(rst), .Q(
        \regs[11][20] ) );
  DFFRHQX1 \regs_reg[11][19]  ( .D(n457), .CK(clk), .RN(rst), .Q(
        \regs[11][19] ) );
  DFFRHQX1 \regs_reg[11][18]  ( .D(n456), .CK(clk), .RN(rst), .Q(
        \regs[11][18] ) );
  DFFRHQX1 \regs_reg[11][17]  ( .D(n455), .CK(clk), .RN(rst), .Q(
        \regs[11][17] ) );
  DFFRHQX1 \regs_reg[11][16]  ( .D(n454), .CK(clk), .RN(rst), .Q(
        \regs[11][16] ) );
  DFFRHQX1 \regs_reg[7][23]  ( .D(n333), .CK(clk), .RN(rst), .Q(\regs[7][23] )
         );
  DFFRHQX1 \regs_reg[7][22]  ( .D(n332), .CK(clk), .RN(rst), .Q(\regs[7][22] )
         );
  DFFRHQX1 \regs_reg[7][21]  ( .D(n331), .CK(clk), .RN(rst), .Q(\regs[7][21] )
         );
  DFFRHQX1 \regs_reg[7][20]  ( .D(n330), .CK(clk), .RN(rst), .Q(\regs[7][20] )
         );
  DFFRHQX1 \regs_reg[7][19]  ( .D(n329), .CK(clk), .RN(rst), .Q(\regs[7][19] )
         );
  DFFRHQX1 \regs_reg[7][18]  ( .D(n328), .CK(clk), .RN(rst), .Q(\regs[7][18] )
         );
  DFFRHQX1 \regs_reg[7][17]  ( .D(n327), .CK(clk), .RN(rst), .Q(\regs[7][17] )
         );
  DFFRHQX1 \regs_reg[7][16]  ( .D(n326), .CK(clk), .RN(rst), .Q(\regs[7][16] )
         );
  DFFRHQX1 \regs_reg[3][23]  ( .D(n205), .CK(clk), .RN(rst), .Q(\regs[3][23] )
         );
  DFFRHQX1 \regs_reg[3][22]  ( .D(n204), .CK(clk), .RN(rst), .Q(\regs[3][22] )
         );
  DFFRHQX1 \regs_reg[3][21]  ( .D(n203), .CK(clk), .RN(rst), .Q(\regs[3][21] )
         );
  DFFRHQX1 \regs_reg[3][20]  ( .D(n202), .CK(clk), .RN(rst), .Q(\regs[3][20] )
         );
  DFFRHQX1 \regs_reg[3][18]  ( .D(n200), .CK(clk), .RN(rst), .Q(\regs[3][18] )
         );
  DFFRHQX1 \regs_reg[3][17]  ( .D(n199), .CK(clk), .RN(rst), .Q(\regs[3][17] )
         );
  DFFRHQX1 \regs_reg[3][16]  ( .D(n198), .CK(clk), .RN(rst), .Q(\regs[3][16] )
         );
  DFFRHQX1 \regs_reg[28][23]  ( .D(n1005), .CK(clk), .RN(rst), .Q(
        \regs[28][23] ) );
  DFFRHQX1 \regs_reg[28][22]  ( .D(n1004), .CK(clk), .RN(rst), .Q(
        \regs[28][22] ) );
  DFFRHQX1 \regs_reg[28][21]  ( .D(n1003), .CK(clk), .RN(rst), .Q(
        \regs[28][21] ) );
  DFFRHQX1 \regs_reg[28][20]  ( .D(n1002), .CK(clk), .RN(rst), .Q(
        \regs[28][20] ) );
  DFFRHQX1 \regs_reg[28][19]  ( .D(n1001), .CK(clk), .RN(rst), .Q(
        \regs[28][19] ) );
  DFFRHQX1 \regs_reg[28][18]  ( .D(n1000), .CK(clk), .RN(rst), .Q(
        \regs[28][18] ) );
  DFFRHQX1 \regs_reg[28][17]  ( .D(n999), .CK(clk), .RN(rst), .Q(
        \regs[28][17] ) );
  DFFRHQX1 \regs_reg[28][16]  ( .D(n998), .CK(clk), .RN(rst), .Q(
        \regs[28][16] ) );
  DFFRHQX1 \regs_reg[24][23]  ( .D(n877), .CK(clk), .RN(rst), .Q(
        \regs[24][23] ) );
  DFFRHQX1 \regs_reg[24][22]  ( .D(n876), .CK(clk), .RN(rst), .Q(
        \regs[24][22] ) );
  DFFRHQX1 \regs_reg[24][21]  ( .D(n875), .CK(clk), .RN(rst), .Q(
        \regs[24][21] ) );
  DFFRHQX1 \regs_reg[24][20]  ( .D(n874), .CK(clk), .RN(rst), .Q(
        \regs[24][20] ) );
  DFFRHQX1 \regs_reg[24][18]  ( .D(n872), .CK(clk), .RN(rst), .Q(
        \regs[24][18] ) );
  DFFRHQX1 \regs_reg[24][17]  ( .D(n871), .CK(clk), .RN(rst), .Q(
        \regs[24][17] ) );
  DFFRHQX1 \regs_reg[24][16]  ( .D(n870), .CK(clk), .RN(rst), .Q(
        \regs[24][16] ) );
  DFFRHQX1 \regs_reg[20][23]  ( .D(n749), .CK(clk), .RN(rst), .Q(
        \regs[20][23] ) );
  DFFRHQX1 \regs_reg[20][22]  ( .D(n748), .CK(clk), .RN(rst), .Q(
        \regs[20][22] ) );
  DFFRHQX1 \regs_reg[20][21]  ( .D(n747), .CK(clk), .RN(rst), .Q(
        \regs[20][21] ) );
  DFFRHQX1 \regs_reg[20][20]  ( .D(n746), .CK(clk), .RN(rst), .Q(
        \regs[20][20] ) );
  DFFRHQX1 \regs_reg[20][19]  ( .D(n745), .CK(clk), .RN(rst), .Q(
        \regs[20][19] ) );
  DFFRHQX1 \regs_reg[20][18]  ( .D(n744), .CK(clk), .RN(rst), .Q(
        \regs[20][18] ) );
  DFFRHQX1 \regs_reg[20][17]  ( .D(n743), .CK(clk), .RN(rst), .Q(
        \regs[20][17] ) );
  DFFRHQX1 \regs_reg[20][16]  ( .D(n742), .CK(clk), .RN(rst), .Q(
        \regs[20][16] ) );
  DFFRHQX1 \regs_reg[16][23]  ( .D(n621), .CK(clk), .RN(rst), .Q(
        \regs[16][23] ) );
  DFFRHQX1 \regs_reg[16][22]  ( .D(n620), .CK(clk), .RN(rst), .Q(
        \regs[16][22] ) );
  DFFRHQX1 \regs_reg[16][21]  ( .D(n619), .CK(clk), .RN(rst), .Q(
        \regs[16][21] ) );
  DFFRHQX1 \regs_reg[16][20]  ( .D(n618), .CK(clk), .RN(rst), .Q(
        \regs[16][20] ) );
  DFFRHQX1 \regs_reg[16][17]  ( .D(n615), .CK(clk), .RN(rst), .Q(
        \regs[16][17] ) );
  DFFRHQX1 \regs_reg[16][16]  ( .D(n614), .CK(clk), .RN(rst), .Q(
        \regs[16][16] ) );
  DFFRHQX1 \regs_reg[12][23]  ( .D(n493), .CK(clk), .RN(rst), .Q(
        \regs[12][23] ) );
  DFFRHQX1 \regs_reg[12][22]  ( .D(n492), .CK(clk), .RN(rst), .Q(
        \regs[12][22] ) );
  DFFRHQX1 \regs_reg[12][21]  ( .D(n491), .CK(clk), .RN(rst), .Q(
        \regs[12][21] ) );
  DFFRHQX1 \regs_reg[12][20]  ( .D(n490), .CK(clk), .RN(rst), .Q(
        \regs[12][20] ) );
  DFFRHQX1 \regs_reg[12][18]  ( .D(n488), .CK(clk), .RN(rst), .Q(
        \regs[12][18] ) );
  DFFRHQX1 \regs_reg[12][17]  ( .D(n487), .CK(clk), .RN(rst), .Q(
        \regs[12][17] ) );
  DFFRHQX1 \regs_reg[12][16]  ( .D(n486), .CK(clk), .RN(rst), .Q(
        \regs[12][16] ) );
  DFFRHQX1 \regs_reg[8][23]  ( .D(n365), .CK(clk), .RN(rst), .Q(\regs[8][23] )
         );
  DFFRHQX1 \regs_reg[8][22]  ( .D(n364), .CK(clk), .RN(rst), .Q(\regs[8][22] )
         );
  DFFRHQX1 \regs_reg[8][21]  ( .D(n363), .CK(clk), .RN(rst), .Q(\regs[8][21] )
         );
  DFFRHQX1 \regs_reg[8][20]  ( .D(n362), .CK(clk), .RN(rst), .Q(\regs[8][20] )
         );
  DFFRHQX1 \regs_reg[8][17]  ( .D(n359), .CK(clk), .RN(rst), .Q(\regs[8][17] )
         );
  DFFRHQX1 \regs_reg[8][16]  ( .D(n358), .CK(clk), .RN(rst), .Q(\regs[8][16] )
         );
  DFFRHQX1 \regs_reg[4][23]  ( .D(n237), .CK(clk), .RN(rst), .Q(\regs[4][23] )
         );
  DFFRHQX1 \regs_reg[4][22]  ( .D(n236), .CK(clk), .RN(rst), .Q(\regs[4][22] )
         );
  DFFRHQX1 \regs_reg[4][21]  ( .D(n235), .CK(clk), .RN(rst), .Q(\regs[4][21] )
         );
  DFFRHQX1 \regs_reg[4][20]  ( .D(n234), .CK(clk), .RN(rst), .Q(\regs[4][20] )
         );
  DFFRHQX1 \regs_reg[4][17]  ( .D(n231), .CK(clk), .RN(rst), .Q(\regs[4][17] )
         );
  DFFRHQX1 \regs_reg[4][16]  ( .D(n230), .CK(clk), .RN(rst), .Q(\regs[4][16] )
         );
  DFFRHQX1 \regs_reg[0][23]  ( .D(n109), .CK(clk), .RN(rst), .Q(\regs[0][23] )
         );
  DFFRHQX1 \regs_reg[0][22]  ( .D(n108), .CK(clk), .RN(rst), .Q(\regs[0][22] )
         );
  DFFRHQX1 \regs_reg[0][21]  ( .D(n107), .CK(clk), .RN(rst), .Q(\regs[0][21] )
         );
  DFFRHQX1 \regs_reg[0][20]  ( .D(n106), .CK(clk), .RN(rst), .Q(\regs[0][20] )
         );
  DFFRHQX1 \regs_reg[30][23]  ( .D(n1069), .CK(clk), .RN(rst), .Q(
        \regs[30][23] ) );
  DFFRHQX1 \regs_reg[30][22]  ( .D(n1068), .CK(clk), .RN(rst), .Q(
        \regs[30][22] ) );
  DFFRHQX1 \regs_reg[30][21]  ( .D(n1067), .CK(clk), .RN(rst), .Q(
        \regs[30][21] ) );
  DFFRHQX1 \regs_reg[30][20]  ( .D(n1066), .CK(clk), .RN(rst), .Q(
        \regs[30][20] ) );
  DFFRHQX1 \regs_reg[30][19]  ( .D(n1065), .CK(clk), .RN(rst), .Q(
        \regs[30][19] ) );
  DFFRHQX1 \regs_reg[30][18]  ( .D(n1064), .CK(clk), .RN(rst), .Q(
        \regs[30][18] ) );
  DFFRHQX1 \regs_reg[30][17]  ( .D(n1063), .CK(clk), .RN(rst), .Q(
        \regs[30][17] ) );
  DFFRHQX1 \regs_reg[30][16]  ( .D(n1062), .CK(clk), .RN(rst), .Q(
        \regs[30][16] ) );
  DFFRHQX1 \regs_reg[26][23]  ( .D(n941), .CK(clk), .RN(rst), .Q(
        \regs[26][23] ) );
  DFFRHQX1 \regs_reg[26][22]  ( .D(n940), .CK(clk), .RN(rst), .Q(
        \regs[26][22] ) );
  DFFRHQX1 \regs_reg[26][21]  ( .D(n939), .CK(clk), .RN(rst), .Q(
        \regs[26][21] ) );
  DFFRHQX1 \regs_reg[26][20]  ( .D(n938), .CK(clk), .RN(rst), .Q(
        \regs[26][20] ) );
  DFFRHQX1 \regs_reg[26][19]  ( .D(n937), .CK(clk), .RN(rst), .Q(
        \regs[26][19] ) );
  DFFRHQX1 \regs_reg[26][18]  ( .D(n936), .CK(clk), .RN(rst), .Q(
        \regs[26][18] ) );
  DFFRHQX1 \regs_reg[26][17]  ( .D(n935), .CK(clk), .RN(rst), .Q(
        \regs[26][17] ) );
  DFFRHQX1 \regs_reg[26][16]  ( .D(n934), .CK(clk), .RN(rst), .Q(
        \regs[26][16] ) );
  DFFRHQX1 \regs_reg[22][23]  ( .D(n813), .CK(clk), .RN(rst), .Q(
        \regs[22][23] ) );
  DFFRHQX1 \regs_reg[22][22]  ( .D(n812), .CK(clk), .RN(rst), .Q(
        \regs[22][22] ) );
  DFFRHQX1 \regs_reg[22][21]  ( .D(n811), .CK(clk), .RN(rst), .Q(
        \regs[22][21] ) );
  DFFRHQX1 \regs_reg[22][20]  ( .D(n810), .CK(clk), .RN(rst), .Q(
        \regs[22][20] ) );
  DFFRHQX1 \regs_reg[22][19]  ( .D(n809), .CK(clk), .RN(rst), .Q(
        \regs[22][19] ) );
  DFFRHQX1 \regs_reg[22][18]  ( .D(n808), .CK(clk), .RN(rst), .Q(
        \regs[22][18] ) );
  DFFRHQX1 \regs_reg[22][17]  ( .D(n807), .CK(clk), .RN(rst), .Q(
        \regs[22][17] ) );
  DFFRHQX1 \regs_reg[22][16]  ( .D(n806), .CK(clk), .RN(rst), .Q(
        \regs[22][16] ) );
  DFFRHQX1 \regs_reg[18][23]  ( .D(n685), .CK(clk), .RN(rst), .Q(
        \regs[18][23] ) );
  DFFRHQX1 \regs_reg[18][22]  ( .D(n684), .CK(clk), .RN(rst), .Q(
        \regs[18][22] ) );
  DFFRHQX1 \regs_reg[18][21]  ( .D(n683), .CK(clk), .RN(rst), .Q(
        \regs[18][21] ) );
  DFFRHQX1 \regs_reg[18][20]  ( .D(n682), .CK(clk), .RN(rst), .Q(
        \regs[18][20] ) );
  DFFRHQX1 \regs_reg[18][19]  ( .D(n681), .CK(clk), .RN(rst), .Q(
        \regs[18][19] ) );
  DFFRHQX1 \regs_reg[18][18]  ( .D(n680), .CK(clk), .RN(rst), .Q(
        \regs[18][18] ) );
  DFFRHQX1 \regs_reg[18][17]  ( .D(n679), .CK(clk), .RN(rst), .Q(
        \regs[18][17] ) );
  DFFRHQX1 \regs_reg[18][16]  ( .D(n678), .CK(clk), .RN(rst), .Q(
        \regs[18][16] ) );
  DFFRHQX1 \regs_reg[14][23]  ( .D(n557), .CK(clk), .RN(rst), .Q(
        \regs[14][23] ) );
  DFFRHQX1 \regs_reg[14][22]  ( .D(n556), .CK(clk), .RN(rst), .Q(
        \regs[14][22] ) );
  DFFRHQX1 \regs_reg[14][21]  ( .D(n555), .CK(clk), .RN(rst), .Q(
        \regs[14][21] ) );
  DFFRHQX1 \regs_reg[14][20]  ( .D(n554), .CK(clk), .RN(rst), .Q(
        \regs[14][20] ) );
  DFFRHQX1 \regs_reg[14][19]  ( .D(n553), .CK(clk), .RN(rst), .Q(
        \regs[14][19] ) );
  DFFRHQX1 \regs_reg[14][18]  ( .D(n552), .CK(clk), .RN(rst), .Q(
        \regs[14][18] ) );
  DFFRHQX1 \regs_reg[14][17]  ( .D(n551), .CK(clk), .RN(rst), .Q(
        \regs[14][17] ) );
  DFFRHQX1 \regs_reg[14][16]  ( .D(n550), .CK(clk), .RN(rst), .Q(
        \regs[14][16] ) );
  DFFRHQX1 \regs_reg[10][23]  ( .D(n429), .CK(clk), .RN(rst), .Q(
        \regs[10][23] ) );
  DFFRHQX1 \regs_reg[10][22]  ( .D(n428), .CK(clk), .RN(rst), .Q(
        \regs[10][22] ) );
  DFFRHQX1 \regs_reg[10][21]  ( .D(n427), .CK(clk), .RN(rst), .Q(
        \regs[10][21] ) );
  DFFRHQX1 \regs_reg[10][20]  ( .D(n426), .CK(clk), .RN(rst), .Q(
        \regs[10][20] ) );
  DFFRHQX1 \regs_reg[10][18]  ( .D(n424), .CK(clk), .RN(rst), .Q(
        \regs[10][18] ) );
  DFFRHQX1 \regs_reg[10][17]  ( .D(n423), .CK(clk), .RN(rst), .Q(
        \regs[10][17] ) );
  DFFRHQX1 \regs_reg[10][16]  ( .D(n422), .CK(clk), .RN(rst), .Q(
        \regs[10][16] ) );
  DFFRHQX1 \regs_reg[6][23]  ( .D(n301), .CK(clk), .RN(rst), .Q(\regs[6][23] )
         );
  DFFRHQX1 \regs_reg[6][22]  ( .D(n300), .CK(clk), .RN(rst), .Q(\regs[6][22] )
         );
  DFFRHQX1 \regs_reg[6][21]  ( .D(n299), .CK(clk), .RN(rst), .Q(\regs[6][21] )
         );
  DFFRHQX1 \regs_reg[6][20]  ( .D(n298), .CK(clk), .RN(rst), .Q(\regs[6][20] )
         );
  DFFRHQX1 \regs_reg[6][19]  ( .D(n297), .CK(clk), .RN(rst), .Q(\regs[6][19] )
         );
  DFFRHQX1 \regs_reg[6][18]  ( .D(n296), .CK(clk), .RN(rst), .Q(\regs[6][18] )
         );
  DFFRHQX1 \regs_reg[6][17]  ( .D(n295), .CK(clk), .RN(rst), .Q(\regs[6][17] )
         );
  DFFRHQX1 \regs_reg[6][16]  ( .D(n294), .CK(clk), .RN(rst), .Q(\regs[6][16] )
         );
  DFFRHQX1 \regs_reg[2][23]  ( .D(n173), .CK(clk), .RN(rst), .Q(\regs[2][23] )
         );
  DFFRHQX1 \regs_reg[2][22]  ( .D(n172), .CK(clk), .RN(rst), .Q(\regs[2][22] )
         );
  DFFRHQX1 \regs_reg[2][21]  ( .D(n171), .CK(clk), .RN(rst), .Q(\regs[2][21] )
         );
  DFFRHQX1 \regs_reg[2][20]  ( .D(n170), .CK(clk), .RN(rst), .Q(\regs[2][20] )
         );
  DFFRHQX1 \regs_reg[2][17]  ( .D(n167), .CK(clk), .RN(rst), .Q(\regs[2][17] )
         );
  DFFRHQX1 \regs_reg[2][16]  ( .D(n166), .CK(clk), .RN(rst), .Q(\regs[2][16] )
         );
  INVXL U2 ( .A(N24), .Y(n2154) );
  INVXL U3 ( .A(N14), .Y(n1409) );
  NAND2X1 U4 ( .A(n38), .B(n36), .Y(n1) );
  NAND2X1 U5 ( .A(n40), .B(n36), .Y(n3) );
  NAND2X1 U6 ( .A(n42), .B(n36), .Y(n4) );
  NAND2X1 U7 ( .A(n46), .B(n35), .Y(n5) );
  NAND2X1 U8 ( .A(n46), .B(n38), .Y(n13) );
  NAND2X1 U9 ( .A(n46), .B(n40), .Y(n14) );
  NAND2X1 U10 ( .A(n46), .B(n42), .Y(n15) );
  NAND2X1 U11 ( .A(n52), .B(n35), .Y(n16) );
  NAND2X1 U12 ( .A(n52), .B(n38), .Y(n17) );
  NAND2X1 U13 ( .A(n52), .B(n40), .Y(n18) );
  NAND2X1 U14 ( .A(n52), .B(n42), .Y(n19) );
  NAND2X1 U15 ( .A(n58), .B(n35), .Y(n20) );
  NAND2X1 U16 ( .A(n58), .B(n38), .Y(n21) );
  NAND2X1 U17 ( .A(n64), .B(n35), .Y(n22) );
  NAND2X1 U18 ( .A(n64), .B(n38), .Y(n23) );
  NAND2X1 U19 ( .A(n58), .B(n40), .Y(n24) );
  NAND2X1 U20 ( .A(n70), .B(n35), .Y(n25) );
  NAND2X1 U21 ( .A(n70), .B(n38), .Y(n26) );
  NAND2X1 U22 ( .A(n70), .B(n40), .Y(n27) );
  NAND2X1 U23 ( .A(n70), .B(n42), .Y(n28) );
  NAND2X1 U24 ( .A(n76), .B(n35), .Y(n29) );
  NAND2X1 U25 ( .A(n76), .B(n38), .Y(n30) );
  NAND2X1 U26 ( .A(n76), .B(n40), .Y(n31) );
  NAND2X1 U27 ( .A(n76), .B(n42), .Y(n32) );
  NAND2X1 U28 ( .A(n81), .B(n35), .Y(n33) );
  NAND2X1 U29 ( .A(n81), .B(n38), .Y(n37) );
  NAND2X1 U30 ( .A(n81), .B(n40), .Y(n39) );
  NAND2X1 U31 ( .A(n81), .B(n42), .Y(n41) );
  INVX1 U32 ( .A(n2181), .Y(n2183) );
  INVX1 U33 ( .A(n2182), .Y(n2184) );
  INVX1 U34 ( .A(n2182), .Y(n2185) );
  INVX1 U35 ( .A(n2182), .Y(n2186) );
  INVX1 U36 ( .A(n2182), .Y(n2187) );
  INVX1 U37 ( .A(n2181), .Y(n2188) );
  INVX1 U38 ( .A(n2181), .Y(n2189) );
  INVX1 U39 ( .A(n2180), .Y(n2190) );
  INVX1 U40 ( .A(n2180), .Y(n2191) );
  INVX1 U41 ( .A(n2180), .Y(n2192) );
  INVX1 U42 ( .A(n2182), .Y(n2193) );
  INVX1 U43 ( .A(n2181), .Y(n2194) );
  INVX1 U44 ( .A(n2181), .Y(n2195) );
  INVX1 U45 ( .A(n2180), .Y(n2196) );
  INVX1 U46 ( .A(n2180), .Y(n2197) );
  INVX1 U47 ( .A(n2181), .Y(n2198) );
  INVX1 U48 ( .A(n2180), .Y(n2199) );
  INVX1 U49 ( .A(n2182), .Y(n2200) );
  INVX1 U50 ( .A(n2182), .Y(n2201) );
  INVX1 U51 ( .A(n2182), .Y(n2202) );
  INVX1 U52 ( .A(n2181), .Y(n2203) );
  INVX1 U53 ( .A(n1437), .Y(n1438) );
  INVX1 U54 ( .A(n1437), .Y(n1439) );
  INVX1 U55 ( .A(n1437), .Y(n1440) );
  INVX1 U56 ( .A(n1437), .Y(n1441) );
  INVX1 U57 ( .A(n1437), .Y(n1442) );
  INVX1 U58 ( .A(n1436), .Y(n1443) );
  INVX1 U59 ( .A(n1437), .Y(n1444) );
  INVX1 U60 ( .A(n1436), .Y(n1445) );
  INVX1 U61 ( .A(n1436), .Y(n1446) );
  INVX1 U62 ( .A(n1436), .Y(n1447) );
  INVX1 U63 ( .A(n1435), .Y(n1448) );
  INVX1 U64 ( .A(n1435), .Y(n1449) );
  INVX1 U65 ( .A(n1435), .Y(n1450) );
  INVX1 U66 ( .A(n1435), .Y(n1451) );
  INVX1 U67 ( .A(n1435), .Y(n1452) );
  INVX1 U68 ( .A(n1435), .Y(n1453) );
  INVX1 U69 ( .A(n1436), .Y(n1454) );
  INVX1 U70 ( .A(n1437), .Y(n1455) );
  INVX1 U71 ( .A(n1436), .Y(n1456) );
  INVX1 U72 ( .A(n1437), .Y(n1457) );
  INVX1 U73 ( .A(n1436), .Y(n1458) );
  INVX1 U74 ( .A(n2157), .Y(n2158) );
  INVX1 U75 ( .A(n2157), .Y(n2159) );
  INVX1 U76 ( .A(n2157), .Y(n2160) );
  INVX1 U77 ( .A(n2157), .Y(n2161) );
  INVX1 U78 ( .A(n2156), .Y(n2162) );
  INVX1 U79 ( .A(n2157), .Y(n2163) );
  INVX1 U80 ( .A(n2157), .Y(n2164) );
  INVX1 U81 ( .A(n2157), .Y(n2165) );
  INVX1 U82 ( .A(n2157), .Y(n2166) );
  INVX1 U83 ( .A(n2157), .Y(n2167) );
  INVX1 U84 ( .A(n2179), .Y(n2168) );
  INVX1 U85 ( .A(n2179), .Y(n2169) );
  INVX1 U86 ( .A(n2179), .Y(n2170) );
  INVX1 U87 ( .A(n2179), .Y(n2171) );
  INVX1 U88 ( .A(n2156), .Y(n2172) );
  INVX1 U89 ( .A(n2179), .Y(n2173) );
  INVX1 U90 ( .A(n2179), .Y(n2174) );
  INVX1 U91 ( .A(n2156), .Y(n2175) );
  INVX1 U92 ( .A(n2156), .Y(n2176) );
  INVX1 U93 ( .A(n2156), .Y(n2177) );
  INVX1 U94 ( .A(n2156), .Y(n2178) );
  INVX1 U95 ( .A(n1413), .Y(n1414) );
  INVX1 U96 ( .A(n1413), .Y(n1415) );
  INVX1 U97 ( .A(n1413), .Y(n1416) );
  INVX1 U98 ( .A(n1413), .Y(n1417) );
  INVX1 U99 ( .A(n1413), .Y(n1418) );
  INVX1 U100 ( .A(n1412), .Y(n1419) );
  INVX1 U101 ( .A(n1412), .Y(n1420) );
  INVX1 U102 ( .A(n1413), .Y(n1421) );
  INVX1 U103 ( .A(n1413), .Y(n1422) );
  INVX1 U104 ( .A(n1412), .Y(n1423) );
  INVX1 U105 ( .A(n1411), .Y(n1424) );
  INVX1 U106 ( .A(n1411), .Y(n1425) );
  INVX1 U107 ( .A(n1411), .Y(n1426) );
  INVX1 U108 ( .A(n1411), .Y(n1427) );
  INVX1 U109 ( .A(n1411), .Y(n1428) );
  INVX1 U110 ( .A(n1411), .Y(n1429) );
  INVX1 U111 ( .A(n1412), .Y(n1430) );
  INVX1 U112 ( .A(n1413), .Y(n1431) );
  INVX1 U113 ( .A(n1412), .Y(n1432) );
  INVX1 U114 ( .A(n1412), .Y(n1433) );
  INVX1 U115 ( .A(n1412), .Y(n1434) );
  INVX1 U116 ( .A(n1807), .Y(n1809) );
  INVX1 U117 ( .A(n1807), .Y(n1810) );
  INVX1 U118 ( .A(n1807), .Y(n1811) );
  INVX1 U119 ( .A(n1807), .Y(n1812) );
  INVX1 U120 ( .A(n1807), .Y(n1813) );
  INVX1 U121 ( .A(n1807), .Y(n1814) );
  INVX1 U122 ( .A(n1807), .Y(n1815) );
  INVX1 U123 ( .A(n1807), .Y(n1816) );
  INVX1 U124 ( .A(n1807), .Y(n1817) );
  INVX1 U125 ( .A(n1807), .Y(n1818) );
  INVX1 U126 ( .A(n1807), .Y(n1819) );
  INVX1 U127 ( .A(n1807), .Y(n1820) );
  INVX1 U128 ( .A(n1807), .Y(n1821) );
  INVX1 U129 ( .A(n1807), .Y(n1822) );
  INVX1 U130 ( .A(n1807), .Y(n1823) );
  INVX1 U131 ( .A(n1807), .Y(n1824) );
  INVX1 U132 ( .A(n1807), .Y(n1825) );
  INVX1 U133 ( .A(n1807), .Y(n1826) );
  INVX1 U134 ( .A(n1807), .Y(n1827) );
  INVX1 U135 ( .A(n1807), .Y(n1828) );
  INVX1 U136 ( .A(n1807), .Y(n1829) );
  INVX1 U137 ( .A(write_data[2]), .Y(n2225) );
  INVX1 U138 ( .A(write_data[13]), .Y(n2221) );
  INVX1 U139 ( .A(write_data[16]), .Y(n2218) );
  INVX1 U140 ( .A(write_data[17]), .Y(n2217) );
  INVX1 U141 ( .A(write_data[18]), .Y(n2216) );
  INVX1 U142 ( .A(write_data[19]), .Y(n2215) );
  INVX1 U143 ( .A(write_data[20]), .Y(n2214) );
  INVX1 U144 ( .A(write_data[21]), .Y(n2213) );
  INVX1 U145 ( .A(write_data[22]), .Y(n2212) );
  INVX1 U146 ( .A(write_data[23]), .Y(n2211) );
  INVX1 U147 ( .A(write_data[24]), .Y(n2210) );
  INVX1 U148 ( .A(write_data[25]), .Y(n2209) );
  INVX1 U149 ( .A(write_data[26]), .Y(n2208) );
  INVX1 U150 ( .A(write_data[27]), .Y(n2207) );
  INVX1 U151 ( .A(write_data[28]), .Y(n2206) );
  INVX1 U152 ( .A(write_data[29]), .Y(n2205) );
  INVX1 U153 ( .A(write_data[30]), .Y(n2204) );
  INVX1 U154 ( .A(n1785), .Y(n1786) );
  INVX1 U155 ( .A(n1784), .Y(n1787) );
  INVX1 U156 ( .A(n1784), .Y(n1788) );
  INVX1 U157 ( .A(n1784), .Y(n1789) );
  INVX1 U158 ( .A(n1784), .Y(n1790) );
  INVX1 U159 ( .A(n1784), .Y(n1791) );
  INVX1 U160 ( .A(n1784), .Y(n1792) );
  INVX1 U161 ( .A(n1785), .Y(n1793) );
  INVX1 U162 ( .A(n1785), .Y(n1794) );
  INVX1 U163 ( .A(n1785), .Y(n1795) );
  INVX1 U164 ( .A(n1785), .Y(n1796) );
  INVX1 U165 ( .A(n1785), .Y(n1797) );
  INVX1 U166 ( .A(n1785), .Y(n1798) );
  INVX1 U167 ( .A(n1784), .Y(n1799) );
  INVX1 U168 ( .A(n1784), .Y(n1800) );
  INVX1 U169 ( .A(n1784), .Y(n1801) );
  INVX1 U170 ( .A(n1784), .Y(n1802) );
  INVX1 U171 ( .A(n1784), .Y(n1803) );
  INVX1 U172 ( .A(n1784), .Y(n1804) );
  INVX1 U173 ( .A(n1784), .Y(n1805) );
  INVX1 U174 ( .A(n1784), .Y(n1806) );
  INVX1 U175 ( .A(n1807), .Y(n1808) );
  INVX1 U176 ( .A(N23), .Y(n2156) );
  INVX1 U177 ( .A(N22), .Y(n2182) );
  INVX1 U178 ( .A(N22), .Y(n2181) );
  INVX1 U179 ( .A(N23), .Y(n2157) );
  INVX1 U180 ( .A(N22), .Y(n2180) );
  INVX1 U181 ( .A(N12), .Y(n1437) );
  INVX1 U182 ( .A(N13), .Y(n1413) );
  INVX1 U183 ( .A(N13), .Y(n1412) );
  INVX1 U184 ( .A(N12), .Y(n1436) );
  INVX1 U185 ( .A(N12), .Y(n1435) );
  INVX1 U186 ( .A(N13), .Y(n1411) );
  INVX1 U187 ( .A(write_data[0]), .Y(n2227) );
  INVX1 U188 ( .A(write_data[1]), .Y(n2226) );
  INVX1 U189 ( .A(write_data[10]), .Y(n2224) );
  INVX1 U190 ( .A(write_data[11]), .Y(n2223) );
  INVX1 U191 ( .A(write_data[12]), .Y(n2222) );
  INVX1 U192 ( .A(write_data[14]), .Y(n2220) );
  INVX1 U193 ( .A(write_data[15]), .Y(n2219) );
  INVX1 U194 ( .A(N17), .Y(n1807) );
  INVX1 U195 ( .A(N18), .Y(n1784) );
  INVX1 U196 ( .A(N18), .Y(n1785) );
  INVX1 U197 ( .A(n2150), .Y(n2152) );
  INVX1 U198 ( .A(n2150), .Y(n2153) );
  INVX1 U199 ( .A(n1405), .Y(n1406) );
  INVX1 U200 ( .A(n1405), .Y(n1407) );
  INVX1 U201 ( .A(n1405), .Y(n1408) );
  INVX1 U202 ( .A(n2154), .Y(n2155) );
  INVX1 U203 ( .A(n1409), .Y(n1410) );
  INVX1 U204 ( .A(n2150), .Y(n2151) );
  INVX1 U205 ( .A(n1779), .Y(n1780) );
  INVX1 U206 ( .A(n1779), .Y(n1781) );
  INVX1 U207 ( .A(n1782), .Y(n1783) );
  INVX1 U208 ( .A(write_data[3]), .Y(n6) );
  INVX1 U209 ( .A(write_data[4]), .Y(n7) );
  INVX1 U210 ( .A(write_data[5]), .Y(n8) );
  INVX1 U211 ( .A(write_data[6]), .Y(n9) );
  INVX1 U212 ( .A(write_data[7]), .Y(n10) );
  INVX1 U213 ( .A(write_data[8]), .Y(n11) );
  INVX1 U214 ( .A(write_data[9]), .Y(n12) );
  INVX1 U215 ( .A(write_data[31]), .Y(n34) );
  INVX1 U216 ( .A(N23), .Y(n2179) );
  INVX1 U217 ( .A(N25), .Y(n2150) );
  INVX1 U218 ( .A(N15), .Y(n1405) );
  INVX1 U219 ( .A(N20), .Y(n1779) );
  INVX1 U220 ( .A(N19), .Y(n1782) );
  AND2X2 U221 ( .A(n50), .B(n43), .Y(n46) );
  AND2X2 U222 ( .A(n56), .B(n43), .Y(n52) );
  AND2X2 U223 ( .A(n62), .B(n43), .Y(n58) );
  AND2X2 U224 ( .A(n68), .B(n44), .Y(n64) );
  AND2X2 U225 ( .A(n68), .B(n50), .Y(n70) );
  AND2X2 U226 ( .A(n68), .B(n56), .Y(n76) );
  AND2X2 U227 ( .A(n68), .B(n62), .Y(n81) );
  AND2X2 U228 ( .A(n43), .B(n44), .Y(n36) );
  NAND2X1 U229 ( .A(n35), .B(n36), .Y(n2) );
  NAND2X1 U230 ( .A(n58), .B(n42), .Y(n61) );
  NAND2X1 U231 ( .A(n64), .B(n42), .Y(n67) );
  NAND2X1 U232 ( .A(n64), .B(n40), .Y(n66) );
  AND2X2 U233 ( .A(N1160), .B(reg_ena), .Y(read_data3[21]) );
  MX2X1 U234 ( .A(n2049), .B(n2044), .S0(N26), .Y(N1160) );
  AND2X2 U235 ( .A(N1159), .B(reg_ena), .Y(read_data3[22]) );
  MX2X1 U236 ( .A(n2059), .B(n2054), .S0(N26), .Y(N1159) );
  AND2X2 U237 ( .A(N1158), .B(reg_ena), .Y(read_data3[23]) );
  MX2X1 U238 ( .A(n2069), .B(n2064), .S0(N26), .Y(N1158) );
  AND2X2 U239 ( .A(N1157), .B(reg_ena), .Y(read_data3[24]) );
  MX2X1 U240 ( .A(n2079), .B(n2074), .S0(N26), .Y(N1157) );
  AND2X2 U241 ( .A(N1156), .B(reg_ena), .Y(read_data3[25]) );
  MX2X1 U242 ( .A(n2089), .B(n2084), .S0(N26), .Y(N1156) );
  AND2X2 U243 ( .A(N1155), .B(reg_ena), .Y(read_data3[26]) );
  MX2X1 U244 ( .A(n2099), .B(n2094), .S0(N26), .Y(N1155) );
  AND2X2 U245 ( .A(N1154), .B(reg_ena), .Y(read_data3[27]) );
  MX2X1 U246 ( .A(n2109), .B(n2104), .S0(N26), .Y(N1154) );
  AND2X2 U247 ( .A(N1153), .B(reg_ena), .Y(read_data3[28]) );
  MX2X1 U248 ( .A(n2119), .B(n2114), .S0(N26), .Y(N1153) );
  AND2X2 U249 ( .A(N1152), .B(reg_ena), .Y(read_data3[29]) );
  MX2X1 U250 ( .A(n2129), .B(n2124), .S0(N26), .Y(N1152) );
  AND2X2 U251 ( .A(N1151), .B(reg_ena), .Y(read_data3[30]) );
  MX2X1 U252 ( .A(n2139), .B(n2134), .S0(N26), .Y(N1151) );
  AND2X2 U253 ( .A(N1150), .B(reg_ena), .Y(read_data3[31]) );
  MX2X1 U254 ( .A(n2149), .B(n2144), .S0(N26), .Y(N1150) );
  AND2X2 U255 ( .A(N1096), .B(reg_ena), .Y(read_data1[21]) );
  MX2X1 U256 ( .A(n1304), .B(n1299), .S0(N16), .Y(N1096) );
  AND2X2 U257 ( .A(N1095), .B(reg_ena), .Y(read_data1[22]) );
  MX2X1 U258 ( .A(n1314), .B(n1309), .S0(N16), .Y(N1095) );
  AND2X2 U259 ( .A(N1094), .B(reg_ena), .Y(read_data1[23]) );
  MX2X1 U260 ( .A(n1324), .B(n1319), .S0(N16), .Y(N1094) );
  AND2X2 U261 ( .A(N1093), .B(reg_ena), .Y(read_data1[24]) );
  MX2X1 U262 ( .A(n1334), .B(n1329), .S0(N16), .Y(N1093) );
  AND2X2 U263 ( .A(N1092), .B(reg_ena), .Y(read_data1[25]) );
  MX2X1 U264 ( .A(n1344), .B(n1339), .S0(N16), .Y(N1092) );
  AND2X2 U265 ( .A(N1091), .B(reg_ena), .Y(read_data1[26]) );
  AND2X2 U266 ( .A(N1090), .B(reg_ena), .Y(read_data1[27]) );
  AND2X2 U267 ( .A(N1089), .B(reg_ena), .Y(read_data1[28]) );
  AND2X2 U268 ( .A(N1088), .B(reg_ena), .Y(read_data1[29]) );
  AND2X2 U269 ( .A(N1087), .B(reg_ena), .Y(read_data1[30]) );
  MX2X1 U270 ( .A(n1394), .B(n1389), .S0(N16), .Y(N1087) );
  AND2X2 U271 ( .A(N1086), .B(reg_ena), .Y(read_data1[31]) );
  MX2X1 U272 ( .A(n1404), .B(n1399), .S0(N16), .Y(N1086) );
  AND2X2 U273 ( .A(N1116), .B(reg_ena), .Y(read_data1[1]) );
  MX2X1 U274 ( .A(n78), .B(n71), .S0(N16), .Y(N1116) );
  AND2X2 U275 ( .A(N1181), .B(reg_ena), .Y(read_data3[0]) );
  MX2X1 U276 ( .A(n1839), .B(n1834), .S0(N26), .Y(N1181) );
  AND2X2 U277 ( .A(N1117), .B(reg_ena), .Y(read_data1[0]) );
  MX2X1 U278 ( .A(n59), .B(n51), .S0(N16), .Y(N1117) );
  AND2X2 U279 ( .A(N1179), .B(reg_ena), .Y(read_data3[2]) );
  MX2X1 U280 ( .A(n1859), .B(n1854), .S0(N26), .Y(N1179) );
  AND2X2 U281 ( .A(N1178), .B(reg_ena), .Y(read_data3[3]) );
  MX2X1 U282 ( .A(n1869), .B(n1864), .S0(N26), .Y(N1178) );
  AND2X2 U283 ( .A(N1177), .B(reg_ena), .Y(read_data3[4]) );
  MX2X1 U284 ( .A(n1879), .B(n1874), .S0(N26), .Y(N1177) );
  AND2X2 U285 ( .A(N1176), .B(reg_ena), .Y(read_data3[5]) );
  MX2X1 U286 ( .A(n1889), .B(n1884), .S0(N26), .Y(N1176) );
  AND2X2 U287 ( .A(N1175), .B(reg_ena), .Y(read_data3[6]) );
  MX2X1 U288 ( .A(n1899), .B(n1894), .S0(N26), .Y(N1175) );
  AND2X2 U289 ( .A(N1174), .B(reg_ena), .Y(read_data3[7]) );
  MX2X1 U290 ( .A(n1909), .B(n1904), .S0(N26), .Y(N1174) );
  AND2X2 U291 ( .A(N1173), .B(reg_ena), .Y(read_data3[8]) );
  MX2X1 U292 ( .A(n1919), .B(n1914), .S0(N26), .Y(N1173) );
  AND2X2 U293 ( .A(reg_ena), .B(N1172), .Y(read_data3[9]) );
  MX2X1 U294 ( .A(n1929), .B(n1924), .S0(N26), .Y(N1172) );
  AND2X2 U295 ( .A(N1171), .B(reg_ena), .Y(read_data3[10]) );
  MX2X1 U296 ( .A(n1939), .B(n1934), .S0(N26), .Y(N1171) );
  AND2X2 U297 ( .A(N1170), .B(reg_ena), .Y(read_data3[11]) );
  MX2X1 U298 ( .A(n1949), .B(n1944), .S0(N26), .Y(N1170) );
  AND2X2 U299 ( .A(N1169), .B(reg_ena), .Y(read_data3[12]) );
  MX2X1 U300 ( .A(n1959), .B(n1954), .S0(N26), .Y(N1169) );
  AND2X2 U301 ( .A(N1168), .B(reg_ena), .Y(read_data3[13]) );
  MX2X1 U302 ( .A(n1969), .B(n1964), .S0(N26), .Y(N1168) );
  AND2X2 U303 ( .A(N1167), .B(reg_ena), .Y(read_data3[14]) );
  MX2X1 U304 ( .A(n1979), .B(n1974), .S0(N26), .Y(N1167) );
  AND2X2 U305 ( .A(N1166), .B(reg_ena), .Y(read_data3[15]) );
  MX2X1 U306 ( .A(n1989), .B(n1984), .S0(N26), .Y(N1166) );
  AND2X2 U307 ( .A(N1165), .B(reg_ena), .Y(read_data3[16]) );
  MX2X1 U308 ( .A(n1999), .B(n1994), .S0(N26), .Y(N1165) );
  AND2X2 U309 ( .A(N1164), .B(reg_ena), .Y(read_data3[17]) );
  MX2X1 U310 ( .A(n2009), .B(n2004), .S0(N26), .Y(N1164) );
  AND2X2 U311 ( .A(N1163), .B(reg_ena), .Y(read_data3[18]) );
  MX2X1 U312 ( .A(n2019), .B(n2014), .S0(N26), .Y(N1163) );
  AND2X2 U313 ( .A(N1162), .B(reg_ena), .Y(read_data3[19]) );
  MX2X1 U314 ( .A(n2029), .B(n2024), .S0(N26), .Y(N1162) );
  AND2X2 U315 ( .A(N1161), .B(reg_ena), .Y(read_data3[20]) );
  MX2X1 U316 ( .A(n2039), .B(n2034), .S0(N26), .Y(N1161) );
  AND2X2 U317 ( .A(N1115), .B(reg_ena), .Y(read_data1[2]) );
  MX2X1 U318 ( .A(n1114), .B(n85), .S0(N16), .Y(N1115) );
  AND2X2 U319 ( .A(N1114), .B(reg_ena), .Y(read_data1[3]) );
  MX2X1 U320 ( .A(n1124), .B(n1119), .S0(N16), .Y(N1114) );
  AND2X2 U321 ( .A(N1113), .B(reg_ena), .Y(read_data1[4]) );
  MX2X1 U322 ( .A(n1134), .B(n1129), .S0(N16), .Y(N1113) );
  AND2X2 U323 ( .A(N1112), .B(reg_ena), .Y(read_data1[5]) );
  MX2X1 U324 ( .A(n1144), .B(n1139), .S0(N16), .Y(N1112) );
  AND2X2 U325 ( .A(N1111), .B(reg_ena), .Y(read_data1[6]) );
  MX2X1 U326 ( .A(n1154), .B(n1149), .S0(N16), .Y(N1111) );
  AND2X2 U327 ( .A(N1110), .B(reg_ena), .Y(read_data1[7]) );
  MX2X1 U328 ( .A(n1164), .B(n1159), .S0(N16), .Y(N1110) );
  AND2X2 U329 ( .A(N1109), .B(reg_ena), .Y(read_data1[8]) );
  MX2X1 U330 ( .A(n1174), .B(n1169), .S0(N16), .Y(N1109) );
  AND2X2 U331 ( .A(N1108), .B(reg_ena), .Y(read_data1[9]) );
  MX2X1 U332 ( .A(n1184), .B(n1179), .S0(N16), .Y(N1108) );
  AND2X2 U333 ( .A(N1107), .B(reg_ena), .Y(read_data1[10]) );
  MX2X1 U334 ( .A(n1194), .B(n1189), .S0(N16), .Y(N1107) );
  AND2X2 U335 ( .A(N1106), .B(reg_ena), .Y(read_data1[11]) );
  MX2X1 U336 ( .A(n1204), .B(n1199), .S0(N16), .Y(N1106) );
  AND2X2 U337 ( .A(N1105), .B(reg_ena), .Y(read_data1[12]) );
  MX2X1 U338 ( .A(n1214), .B(n1209), .S0(N16), .Y(N1105) );
  AND2X2 U339 ( .A(N1104), .B(reg_ena), .Y(read_data1[13]) );
  MX2X1 U340 ( .A(n1224), .B(n1219), .S0(N16), .Y(N1104) );
  AND2X2 U341 ( .A(N1103), .B(reg_ena), .Y(read_data1[14]) );
  MX2X1 U342 ( .A(n1234), .B(n1229), .S0(N16), .Y(N1103) );
  AND2X2 U343 ( .A(N1102), .B(reg_ena), .Y(read_data1[15]) );
  MX2X1 U344 ( .A(n1244), .B(n1239), .S0(N16), .Y(N1102) );
  AND2X2 U345 ( .A(N1101), .B(reg_ena), .Y(read_data1[16]) );
  MX2X1 U346 ( .A(n1254), .B(n1249), .S0(N16), .Y(N1101) );
  AND2X2 U347 ( .A(N1100), .B(reg_ena), .Y(read_data1[17]) );
  MX2X1 U348 ( .A(n1264), .B(n1259), .S0(N16), .Y(N1100) );
  AND2X2 U349 ( .A(N1099), .B(reg_ena), .Y(read_data1[18]) );
  MX2X1 U350 ( .A(n1274), .B(n1269), .S0(N16), .Y(N1099) );
  AND2X2 U351 ( .A(N1098), .B(reg_ena), .Y(read_data1[19]) );
  MX2X1 U352 ( .A(n1284), .B(n1279), .S0(N16), .Y(N1098) );
  AND2X2 U353 ( .A(N1097), .B(reg_ena), .Y(read_data1[20]) );
  MX2X1 U354 ( .A(n1294), .B(n1289), .S0(N16), .Y(N1097) );
  AND2X2 U355 ( .A(N1180), .B(reg_ena), .Y(read_data3[1]) );
  MX2X1 U356 ( .A(n1849), .B(n1844), .S0(N26), .Y(N1180) );
  MX4X1 U357 ( .A(n1838), .B(n1836), .C(n1837), .D(n1835), .S0(n2151), .S1(
        n2155), .Y(n1839) );
  MX4X1 U358 ( .A(\regs[0][0] ), .B(\regs[1][0] ), .C(\regs[2][0] ), .D(
        \regs[3][0] ), .S0(n2183), .S1(n2158), .Y(n1838) );
  MX4X1 U359 ( .A(\regs[8][0] ), .B(\regs[9][0] ), .C(\regs[10][0] ), .D(
        \regs[11][0] ), .S0(n2183), .S1(n2158), .Y(n1836) );
  MX4X1 U360 ( .A(\regs[4][0] ), .B(\regs[5][0] ), .C(\regs[6][0] ), .D(
        \regs[7][0] ), .S0(n2183), .S1(n2158), .Y(n1837) );
  MX4X1 U361 ( .A(n1848), .B(n1846), .C(n1847), .D(n1845), .S0(n2151), .S1(
        n2155), .Y(n1849) );
  MX4X1 U362 ( .A(\regs[0][1] ), .B(\regs[1][1] ), .C(\regs[2][1] ), .D(
        \regs[3][1] ), .S0(n2183), .S1(n2158), .Y(n1848) );
  MX4X1 U363 ( .A(\regs[8][1] ), .B(\regs[9][1] ), .C(\regs[10][1] ), .D(
        \regs[11][1] ), .S0(n2183), .S1(n2158), .Y(n1846) );
  MX4X1 U364 ( .A(\regs[4][1] ), .B(\regs[5][1] ), .C(\regs[6][1] ), .D(
        \regs[7][1] ), .S0(n2183), .S1(n2158), .Y(n1847) );
  MX4X1 U365 ( .A(n1858), .B(n1856), .C(n1857), .D(n1855), .S0(n2152), .S1(
        n2155), .Y(n1859) );
  MX4X1 U366 ( .A(\regs[0][2] ), .B(\regs[1][2] ), .C(\regs[2][2] ), .D(
        \regs[3][2] ), .S0(n2184), .S1(n2159), .Y(n1858) );
  MX4X1 U367 ( .A(\regs[8][2] ), .B(\regs[9][2] ), .C(\regs[10][2] ), .D(
        \regs[11][2] ), .S0(n2184), .S1(n2159), .Y(n1856) );
  MX4X1 U368 ( .A(\regs[4][2] ), .B(\regs[5][2] ), .C(\regs[6][2] ), .D(
        \regs[7][2] ), .S0(n2184), .S1(n2159), .Y(n1857) );
  MX4X1 U369 ( .A(n1868), .B(n1866), .C(n1867), .D(n1865), .S0(n2152), .S1(
        n2155), .Y(n1869) );
  MX4X1 U370 ( .A(\regs[0][3] ), .B(\regs[1][3] ), .C(\regs[2][3] ), .D(
        \regs[3][3] ), .S0(n2185), .S1(n2160), .Y(n1868) );
  MX4X1 U371 ( .A(\regs[8][3] ), .B(\regs[9][3] ), .C(\regs[10][3] ), .D(
        \regs[11][3] ), .S0(n2185), .S1(n2160), .Y(n1866) );
  MX4X1 U372 ( .A(\regs[4][3] ), .B(\regs[5][3] ), .C(\regs[6][3] ), .D(
        \regs[7][3] ), .S0(n2185), .S1(n2160), .Y(n1867) );
  MX4X1 U373 ( .A(n1878), .B(n1876), .C(n1877), .D(n1875), .S0(n2152), .S1(
        n2155), .Y(n1879) );
  MX4X1 U374 ( .A(\regs[0][4] ), .B(\regs[1][4] ), .C(\regs[2][4] ), .D(
        \regs[3][4] ), .S0(n2185), .S1(n2160), .Y(n1878) );
  MX4X1 U375 ( .A(\regs[8][4] ), .B(\regs[9][4] ), .C(\regs[10][4] ), .D(
        \regs[11][4] ), .S0(n2185), .S1(n2160), .Y(n1876) );
  MX4X1 U376 ( .A(\regs[4][4] ), .B(\regs[5][4] ), .C(\regs[6][4] ), .D(
        \regs[7][4] ), .S0(n2185), .S1(n2160), .Y(n1877) );
  MX4X1 U377 ( .A(n1888), .B(n1886), .C(n1887), .D(n1885), .S0(n2152), .S1(
        n2155), .Y(n1889) );
  MX4X1 U378 ( .A(\regs[0][5] ), .B(\regs[1][5] ), .C(\regs[2][5] ), .D(
        \regs[3][5] ), .S0(n2186), .S1(n2161), .Y(n1888) );
  MX4X1 U379 ( .A(\regs[8][5] ), .B(\regs[9][5] ), .C(\regs[10][5] ), .D(
        \regs[11][5] ), .S0(n2186), .S1(n2161), .Y(n1886) );
  MX4X1 U380 ( .A(\regs[4][5] ), .B(\regs[5][5] ), .C(\regs[6][5] ), .D(
        \regs[7][5] ), .S0(n2186), .S1(n2161), .Y(n1887) );
  MX4X1 U381 ( .A(n1898), .B(n1896), .C(n1897), .D(n1895), .S0(n2152), .S1(
        n2155), .Y(n1899) );
  MX4X1 U382 ( .A(\regs[0][6] ), .B(\regs[1][6] ), .C(\regs[2][6] ), .D(
        \regs[3][6] ), .S0(n2187), .S1(n2162), .Y(n1898) );
  MX4X1 U383 ( .A(\regs[8][6] ), .B(\regs[9][6] ), .C(\regs[10][6] ), .D(
        \regs[11][6] ), .S0(n2187), .S1(n2162), .Y(n1896) );
  MX4X1 U384 ( .A(\regs[4][6] ), .B(\regs[5][6] ), .C(\regs[6][6] ), .D(
        \regs[7][6] ), .S0(n2187), .S1(n2162), .Y(n1897) );
  MX4X1 U385 ( .A(n1908), .B(n1906), .C(n1907), .D(n1905), .S0(n2152), .S1(
        n2155), .Y(n1909) );
  MX4X1 U386 ( .A(\regs[0][7] ), .B(\regs[1][7] ), .C(\regs[2][7] ), .D(
        \regs[3][7] ), .S0(n2187), .S1(n2162), .Y(n1908) );
  MX4X1 U387 ( .A(\regs[8][7] ), .B(\regs[9][7] ), .C(\regs[10][7] ), .D(
        \regs[11][7] ), .S0(n2187), .S1(n2162), .Y(n1906) );
  MX4X1 U388 ( .A(\regs[4][7] ), .B(\regs[5][7] ), .C(\regs[6][7] ), .D(
        \regs[7][7] ), .S0(n2187), .S1(n2162), .Y(n1907) );
  MX4X1 U389 ( .A(n1918), .B(n1916), .C(n1917), .D(n1915), .S0(n2153), .S1(
        n2155), .Y(n1919) );
  MX4X1 U390 ( .A(\regs[0][8] ), .B(\regs[1][8] ), .C(\regs[2][8] ), .D(
        \regs[3][8] ), .S0(n2188), .S1(n2163), .Y(n1918) );
  MX4X1 U391 ( .A(\regs[8][8] ), .B(\regs[9][8] ), .C(\regs[10][8] ), .D(
        \regs[11][8] ), .S0(n2188), .S1(n2163), .Y(n1916) );
  MX4X1 U392 ( .A(\regs[4][8] ), .B(\regs[5][8] ), .C(\regs[6][8] ), .D(
        \regs[7][8] ), .S0(n2188), .S1(n2163), .Y(n1917) );
  MX4X1 U393 ( .A(n1928), .B(n1926), .C(n1927), .D(n1925), .S0(N25), .S1(n2155), .Y(n1929) );
  MX4X1 U394 ( .A(\regs[0][9] ), .B(\regs[1][9] ), .C(\regs[2][9] ), .D(
        \regs[3][9] ), .S0(n2189), .S1(n2164), .Y(n1928) );
  MX4X1 U395 ( .A(\regs[8][9] ), .B(\regs[9][9] ), .C(\regs[10][9] ), .D(
        \regs[11][9] ), .S0(n2189), .S1(n2164), .Y(n1926) );
  MX4X1 U396 ( .A(\regs[4][9] ), .B(\regs[5][9] ), .C(\regs[6][9] ), .D(
        \regs[7][9] ), .S0(n2189), .S1(n2164), .Y(n1927) );
  MX4X1 U397 ( .A(n1938), .B(n1936), .C(n1937), .D(n1935), .S0(N25), .S1(n2155), .Y(n1939) );
  MX4X1 U398 ( .A(\regs[0][10] ), .B(\regs[1][10] ), .C(\regs[2][10] ), .D(
        \regs[3][10] ), .S0(n2189), .S1(n2164), .Y(n1938) );
  MX4X1 U399 ( .A(\regs[8][10] ), .B(\regs[9][10] ), .C(\regs[10][10] ), .D(
        \regs[11][10] ), .S0(n2189), .S1(n2164), .Y(n1936) );
  MX4X1 U400 ( .A(\regs[4][10] ), .B(\regs[5][10] ), .C(\regs[6][10] ), .D(
        \regs[7][10] ), .S0(n2189), .S1(n2164), .Y(n1937) );
  MX4X1 U401 ( .A(n1948), .B(n1946), .C(n1947), .D(n1945), .S0(N25), .S1(n2155), .Y(n1949) );
  MX4X1 U402 ( .A(\regs[0][11] ), .B(\regs[1][11] ), .C(\regs[2][11] ), .D(
        \regs[3][11] ), .S0(n2190), .S1(n2165), .Y(n1948) );
  MX4X1 U403 ( .A(\regs[8][11] ), .B(\regs[9][11] ), .C(\regs[10][11] ), .D(
        \regs[11][11] ), .S0(n2190), .S1(n2165), .Y(n1946) );
  MX4X1 U404 ( .A(\regs[4][11] ), .B(\regs[5][11] ), .C(\regs[6][11] ), .D(
        \regs[7][11] ), .S0(n2190), .S1(n2165), .Y(n1947) );
  MX4X1 U405 ( .A(n1958), .B(n1956), .C(n1957), .D(n1955), .S0(N25), .S1(n2155), .Y(n1959) );
  MX4X1 U406 ( .A(\regs[0][12] ), .B(\regs[1][12] ), .C(\regs[2][12] ), .D(
        \regs[3][12] ), .S0(n2191), .S1(n2166), .Y(n1958) );
  MX4X1 U407 ( .A(\regs[8][12] ), .B(\regs[9][12] ), .C(\regs[10][12] ), .D(
        \regs[11][12] ), .S0(n2191), .S1(n2166), .Y(n1956) );
  MX4X1 U408 ( .A(\regs[4][12] ), .B(\regs[5][12] ), .C(\regs[6][12] ), .D(
        \regs[7][12] ), .S0(n2191), .S1(n2166), .Y(n1957) );
  MX4X1 U409 ( .A(n1968), .B(n1966), .C(n1967), .D(n1965), .S0(n2151), .S1(
        n2155), .Y(n1969) );
  MX4X1 U410 ( .A(\regs[0][13] ), .B(\regs[1][13] ), .C(\regs[2][13] ), .D(
        \regs[3][13] ), .S0(n2191), .S1(n2166), .Y(n1968) );
  MX4X1 U411 ( .A(\regs[8][13] ), .B(\regs[9][13] ), .C(\regs[10][13] ), .D(
        \regs[11][13] ), .S0(n2191), .S1(n2166), .Y(n1966) );
  MX4X1 U412 ( .A(\regs[4][13] ), .B(\regs[5][13] ), .C(\regs[6][13] ), .D(
        \regs[7][13] ), .S0(n2191), .S1(n2166), .Y(n1967) );
  MX4X1 U413 ( .A(n1978), .B(n1976), .C(n1977), .D(n1975), .S0(n2153), .S1(N24), .Y(n1979) );
  MX4X1 U414 ( .A(\regs[0][14] ), .B(\regs[1][14] ), .C(\regs[2][14] ), .D(
        \regs[3][14] ), .S0(n2192), .S1(n2167), .Y(n1978) );
  MX4X1 U415 ( .A(\regs[8][14] ), .B(\regs[9][14] ), .C(\regs[10][14] ), .D(
        \regs[11][14] ), .S0(n2192), .S1(n2167), .Y(n1976) );
  MX4X1 U416 ( .A(\regs[4][14] ), .B(\regs[5][14] ), .C(\regs[6][14] ), .D(
        \regs[7][14] ), .S0(n2192), .S1(n2167), .Y(n1977) );
  MX4X1 U417 ( .A(n1988), .B(n1986), .C(n1987), .D(n1985), .S0(n2153), .S1(N24), .Y(n1989) );
  MX4X1 U418 ( .A(\regs[0][15] ), .B(\regs[1][15] ), .C(\regs[2][15] ), .D(
        \regs[3][15] ), .S0(n2193), .S1(n2168), .Y(n1988) );
  MX4X1 U419 ( .A(\regs[8][15] ), .B(\regs[9][15] ), .C(\regs[10][15] ), .D(
        \regs[11][15] ), .S0(n2193), .S1(n2168), .Y(n1986) );
  MX4X1 U420 ( .A(\regs[4][15] ), .B(\regs[5][15] ), .C(\regs[6][15] ), .D(
        \regs[7][15] ), .S0(n2193), .S1(n2168), .Y(n1987) );
  MX4X1 U421 ( .A(n1998), .B(n1996), .C(n1997), .D(n1995), .S0(n2153), .S1(N24), .Y(n1999) );
  MX4X1 U422 ( .A(\regs[0][16] ), .B(\regs[1][16] ), .C(\regs[2][16] ), .D(
        \regs[3][16] ), .S0(n2193), .S1(n2168), .Y(n1998) );
  MX4X1 U423 ( .A(\regs[8][16] ), .B(\regs[9][16] ), .C(\regs[10][16] ), .D(
        \regs[11][16] ), .S0(n2193), .S1(n2168), .Y(n1996) );
  MX4X1 U424 ( .A(\regs[4][16] ), .B(\regs[5][16] ), .C(\regs[6][16] ), .D(
        \regs[7][16] ), .S0(n2193), .S1(n2168), .Y(n1997) );
  MX4X1 U425 ( .A(n2008), .B(n2006), .C(n2007), .D(n2005), .S0(n2153), .S1(
        n2155), .Y(n2009) );
  MX4X1 U426 ( .A(\regs[0][17] ), .B(\regs[1][17] ), .C(\regs[2][17] ), .D(
        \regs[3][17] ), .S0(n2194), .S1(n2169), .Y(n2008) );
  MX4X1 U427 ( .A(\regs[8][17] ), .B(\regs[9][17] ), .C(\regs[10][17] ), .D(
        \regs[11][17] ), .S0(n2194), .S1(n2169), .Y(n2006) );
  MX4X1 U428 ( .A(\regs[4][17] ), .B(\regs[5][17] ), .C(\regs[6][17] ), .D(
        \regs[7][17] ), .S0(n2194), .S1(n2169), .Y(n2007) );
  MX4X1 U429 ( .A(n2018), .B(n2016), .C(n2017), .D(n2015), .S0(n2153), .S1(N24), .Y(n2019) );
  MX4X1 U430 ( .A(\regs[0][18] ), .B(\regs[1][18] ), .C(\regs[2][18] ), .D(
        \regs[3][18] ), .S0(n2195), .S1(n2170), .Y(n2018) );
  MX4X1 U431 ( .A(\regs[8][18] ), .B(\regs[9][18] ), .C(\regs[10][18] ), .D(
        \regs[11][18] ), .S0(n2195), .S1(n2170), .Y(n2016) );
  MX4X1 U432 ( .A(\regs[4][18] ), .B(\regs[5][18] ), .C(\regs[6][18] ), .D(
        \regs[7][18] ), .S0(n2195), .S1(n2170), .Y(n2017) );
  MX4X1 U433 ( .A(n2028), .B(n2026), .C(n2027), .D(n2025), .S0(n2153), .S1(N24), .Y(n2029) );
  MX4X1 U434 ( .A(\regs[0][19] ), .B(\regs[1][19] ), .C(\regs[2][19] ), .D(
        \regs[3][19] ), .S0(n2195), .S1(n2170), .Y(n2028) );
  MX4X1 U435 ( .A(\regs[8][19] ), .B(\regs[9][19] ), .C(\regs[10][19] ), .D(
        \regs[11][19] ), .S0(n2195), .S1(n2170), .Y(n2026) );
  MX4X1 U436 ( .A(\regs[4][19] ), .B(\regs[5][19] ), .C(\regs[6][19] ), .D(
        \regs[7][19] ), .S0(n2195), .S1(n2170), .Y(n2027) );
  MX4X1 U437 ( .A(n2038), .B(n2036), .C(n2037), .D(n2035), .S0(N25), .S1(N24), 
        .Y(n2039) );
  MX4X1 U438 ( .A(\regs[0][20] ), .B(\regs[1][20] ), .C(\regs[2][20] ), .D(
        \regs[3][20] ), .S0(n2196), .S1(n2171), .Y(n2038) );
  MX4X1 U439 ( .A(\regs[8][20] ), .B(\regs[9][20] ), .C(\regs[10][20] ), .D(
        \regs[11][20] ), .S0(n2196), .S1(n2171), .Y(n2036) );
  MX4X1 U440 ( .A(\regs[4][20] ), .B(\regs[5][20] ), .C(\regs[6][20] ), .D(
        \regs[7][20] ), .S0(n2196), .S1(n2171), .Y(n2037) );
  MX4X1 U441 ( .A(n2048), .B(n2046), .C(n2047), .D(n2045), .S0(N25), .S1(N24), 
        .Y(n2049) );
  MX4X1 U442 ( .A(\regs[0][21] ), .B(\regs[1][21] ), .C(\regs[2][21] ), .D(
        \regs[3][21] ), .S0(n2197), .S1(n2172), .Y(n2048) );
  MX4X1 U443 ( .A(\regs[8][21] ), .B(\regs[9][21] ), .C(\regs[10][21] ), .D(
        \regs[11][21] ), .S0(n2197), .S1(n2172), .Y(n2046) );
  MX4X1 U444 ( .A(\regs[4][21] ), .B(\regs[5][21] ), .C(\regs[6][21] ), .D(
        \regs[7][21] ), .S0(n2197), .S1(n2172), .Y(n2047) );
  MX4X1 U445 ( .A(n2058), .B(n2056), .C(n2057), .D(n2055), .S0(n2151), .S1(N24), .Y(n2059) );
  MX4X1 U446 ( .A(\regs[0][22] ), .B(\regs[1][22] ), .C(\regs[2][22] ), .D(
        \regs[3][22] ), .S0(n2197), .S1(n2172), .Y(n2058) );
  MX4X1 U447 ( .A(\regs[8][22] ), .B(\regs[9][22] ), .C(\regs[10][22] ), .D(
        \regs[11][22] ), .S0(n2197), .S1(n2172), .Y(n2056) );
  MX4X1 U448 ( .A(\regs[4][22] ), .B(\regs[5][22] ), .C(\regs[6][22] ), .D(
        \regs[7][22] ), .S0(n2197), .S1(n2172), .Y(n2057) );
  MX4X1 U449 ( .A(n2068), .B(n2066), .C(n2067), .D(n2065), .S0(N25), .S1(n2155), .Y(n2069) );
  MX4X1 U450 ( .A(\regs[0][23] ), .B(\regs[1][23] ), .C(\regs[2][23] ), .D(
        \regs[3][23] ), .S0(n2198), .S1(n2173), .Y(n2068) );
  MX4X1 U451 ( .A(\regs[8][23] ), .B(\regs[9][23] ), .C(\regs[10][23] ), .D(
        \regs[11][23] ), .S0(n2198), .S1(n2173), .Y(n2066) );
  MX4X1 U452 ( .A(\regs[4][23] ), .B(\regs[5][23] ), .C(\regs[6][23] ), .D(
        \regs[7][23] ), .S0(n2198), .S1(n2173), .Y(n2067) );
  MX4X1 U453 ( .A(n2078), .B(n2076), .C(n2077), .D(n2075), .S0(n2153), .S1(N24), .Y(n2079) );
  MX4X1 U454 ( .A(\regs[0][24] ), .B(\regs[1][24] ), .C(\regs[2][24] ), .D(
        \regs[3][24] ), .S0(n2199), .S1(n2174), .Y(n2078) );
  MX4X1 U455 ( .A(\regs[8][24] ), .B(\regs[9][24] ), .C(\regs[10][24] ), .D(
        \regs[11][24] ), .S0(n2199), .S1(n2174), .Y(n2076) );
  MX4X1 U456 ( .A(\regs[4][24] ), .B(\regs[5][24] ), .C(\regs[6][24] ), .D(
        \regs[7][24] ), .S0(n2199), .S1(n2174), .Y(n2077) );
  MX4X1 U457 ( .A(n2088), .B(n2086), .C(n2087), .D(n2085), .S0(N25), .S1(N24), 
        .Y(n2089) );
  MX4X1 U458 ( .A(\regs[0][25] ), .B(\regs[1][25] ), .C(\regs[2][25] ), .D(
        \regs[3][25] ), .S0(n2199), .S1(n2174), .Y(n2088) );
  MX4X1 U459 ( .A(\regs[8][25] ), .B(\regs[9][25] ), .C(\regs[10][25] ), .D(
        \regs[11][25] ), .S0(n2199), .S1(n2174), .Y(n2086) );
  MX4X1 U460 ( .A(\regs[4][25] ), .B(\regs[5][25] ), .C(\regs[6][25] ), .D(
        \regs[7][25] ), .S0(n2199), .S1(n2174), .Y(n2087) );
  MX4X1 U461 ( .A(n2098), .B(n2096), .C(n2097), .D(n2095), .S0(n2152), .S1(N24), .Y(n2099) );
  MX4X1 U462 ( .A(\regs[0][26] ), .B(\regs[1][26] ), .C(\regs[2][26] ), .D(
        \regs[3][26] ), .S0(n2200), .S1(n2175), .Y(n2098) );
  MX4X1 U463 ( .A(\regs[8][26] ), .B(\regs[9][26] ), .C(\regs[10][26] ), .D(
        \regs[11][26] ), .S0(n2200), .S1(n2175), .Y(n2096) );
  MX4X1 U464 ( .A(\regs[4][26] ), .B(\regs[5][26] ), .C(\regs[6][26] ), .D(
        \regs[7][26] ), .S0(n2200), .S1(n2175), .Y(n2097) );
  MX4X1 U465 ( .A(n2108), .B(n2106), .C(n2107), .D(n2105), .S0(n2152), .S1(
        n2155), .Y(n2109) );
  MX4X1 U466 ( .A(\regs[0][27] ), .B(\regs[1][27] ), .C(\regs[2][27] ), .D(
        \regs[3][27] ), .S0(n2201), .S1(n2176), .Y(n2108) );
  MX4X1 U467 ( .A(\regs[8][27] ), .B(\regs[9][27] ), .C(\regs[10][27] ), .D(
        \regs[11][27] ), .S0(n2201), .S1(n2176), .Y(n2106) );
  MX4X1 U468 ( .A(\regs[4][27] ), .B(\regs[5][27] ), .C(\regs[6][27] ), .D(
        \regs[7][27] ), .S0(n2201), .S1(n2176), .Y(n2107) );
  MX4X1 U469 ( .A(n2118), .B(n2116), .C(n2117), .D(n2115), .S0(n2151), .S1(
        n2155), .Y(n2119) );
  MX4X1 U470 ( .A(\regs[0][28] ), .B(\regs[1][28] ), .C(\regs[2][28] ), .D(
        \regs[3][28] ), .S0(n2201), .S1(n2176), .Y(n2118) );
  MX4X1 U471 ( .A(\regs[8][28] ), .B(\regs[9][28] ), .C(\regs[10][28] ), .D(
        \regs[11][28] ), .S0(n2201), .S1(n2176), .Y(n2116) );
  MX4X1 U472 ( .A(\regs[4][28] ), .B(\regs[5][28] ), .C(\regs[6][28] ), .D(
        \regs[7][28] ), .S0(n2201), .S1(n2176), .Y(n2117) );
  MX4X1 U473 ( .A(n2128), .B(n2126), .C(n2127), .D(n2125), .S0(n2151), .S1(N24), .Y(n2129) );
  MX4X1 U474 ( .A(\regs[0][29] ), .B(\regs[1][29] ), .C(\regs[2][29] ), .D(
        \regs[3][29] ), .S0(n2202), .S1(n2177), .Y(n2128) );
  MX4X1 U475 ( .A(\regs[8][29] ), .B(\regs[9][29] ), .C(\regs[10][29] ), .D(
        \regs[11][29] ), .S0(n2202), .S1(n2177), .Y(n2126) );
  MX4X1 U476 ( .A(\regs[4][29] ), .B(\regs[5][29] ), .C(\regs[6][29] ), .D(
        \regs[7][29] ), .S0(n2202), .S1(n2177), .Y(n2127) );
  MX4X1 U477 ( .A(n2138), .B(n2136), .C(n2137), .D(n2135), .S0(n2151), .S1(N24), .Y(n2139) );
  MX4X1 U478 ( .A(\regs[0][30] ), .B(\regs[1][30] ), .C(\regs[2][30] ), .D(
        \regs[3][30] ), .S0(n2203), .S1(n2178), .Y(n2138) );
  MX4X1 U479 ( .A(\regs[8][30] ), .B(\regs[9][30] ), .C(\regs[10][30] ), .D(
        \regs[11][30] ), .S0(n2203), .S1(n2178), .Y(n2136) );
  MX4X1 U480 ( .A(\regs[4][30] ), .B(\regs[5][30] ), .C(\regs[6][30] ), .D(
        \regs[7][30] ), .S0(n2203), .S1(n2178), .Y(n2137) );
  MX4X1 U481 ( .A(n2148), .B(n2146), .C(n2147), .D(n2145), .S0(n2151), .S1(N24), .Y(n2149) );
  MX4X1 U482 ( .A(\regs[0][31] ), .B(\regs[1][31] ), .C(\regs[2][31] ), .D(
        \regs[3][31] ), .S0(n2203), .S1(n2178), .Y(n2148) );
  MX4X1 U483 ( .A(\regs[8][31] ), .B(\regs[9][31] ), .C(\regs[10][31] ), .D(
        \regs[11][31] ), .S0(n2203), .S1(n2178), .Y(n2146) );
  MX4X1 U484 ( .A(\regs[4][31] ), .B(\regs[5][31] ), .C(\regs[6][31] ), .D(
        \regs[7][31] ), .S0(n2203), .S1(n2178), .Y(n2147) );
  MX4X1 U485 ( .A(n57), .B(n54), .C(n55), .D(n53), .S0(n1406), .S1(n1410), .Y(
        n59) );
  MX4X1 U486 ( .A(\regs[0][0] ), .B(\regs[1][0] ), .C(\regs[2][0] ), .D(
        \regs[3][0] ), .S0(n1438), .S1(n1414), .Y(n57) );
  MX4X1 U487 ( .A(\regs[8][0] ), .B(\regs[9][0] ), .C(\regs[10][0] ), .D(
        \regs[11][0] ), .S0(n1438), .S1(n1414), .Y(n54) );
  MX4X1 U488 ( .A(\regs[4][0] ), .B(\regs[5][0] ), .C(\regs[6][0] ), .D(
        \regs[7][0] ), .S0(n1438), .S1(n1414), .Y(n55) );
  MX4X1 U489 ( .A(n77), .B(n73), .C(n75), .D(n72), .S0(n1406), .S1(n1410), .Y(
        n78) );
  MX4X1 U490 ( .A(\regs[0][1] ), .B(\regs[1][1] ), .C(\regs[2][1] ), .D(
        \regs[3][1] ), .S0(n1438), .S1(n1414), .Y(n77) );
  MX4X1 U491 ( .A(\regs[8][1] ), .B(\regs[9][1] ), .C(\regs[10][1] ), .D(
        \regs[11][1] ), .S0(n1438), .S1(n1414), .Y(n73) );
  MX4X1 U492 ( .A(\regs[4][1] ), .B(\regs[5][1] ), .C(\regs[6][1] ), .D(
        \regs[7][1] ), .S0(n1438), .S1(n1414), .Y(n75) );
  MX4X1 U493 ( .A(n1113), .B(n1111), .C(n1112), .D(n1110), .S0(n1406), .S1(
        n1410), .Y(n1114) );
  MX4X1 U494 ( .A(\regs[0][2] ), .B(\regs[1][2] ), .C(\regs[2][2] ), .D(
        \regs[3][2] ), .S0(n1439), .S1(n1415), .Y(n1113) );
  MX4X1 U495 ( .A(\regs[8][2] ), .B(\regs[9][2] ), .C(\regs[10][2] ), .D(
        \regs[11][2] ), .S0(n1439), .S1(n1415), .Y(n1111) );
  MX4X1 U496 ( .A(\regs[4][2] ), .B(\regs[5][2] ), .C(\regs[6][2] ), .D(
        \regs[7][2] ), .S0(n1439), .S1(n1415), .Y(n1112) );
  MX4X1 U497 ( .A(n1123), .B(n1121), .C(n1122), .D(n1120), .S0(n1406), .S1(
        n1410), .Y(n1124) );
  MX4X1 U498 ( .A(\regs[0][3] ), .B(\regs[1][3] ), .C(\regs[2][3] ), .D(
        \regs[3][3] ), .S0(n1440), .S1(n1416), .Y(n1123) );
  MX4X1 U499 ( .A(\regs[8][3] ), .B(\regs[9][3] ), .C(\regs[10][3] ), .D(
        \regs[11][3] ), .S0(n1440), .S1(n1416), .Y(n1121) );
  MX4X1 U500 ( .A(\regs[4][3] ), .B(\regs[5][3] ), .C(\regs[6][3] ), .D(
        \regs[7][3] ), .S0(n1440), .S1(n1416), .Y(n1122) );
  MX4X1 U501 ( .A(n1133), .B(n1131), .C(n1132), .D(n1130), .S0(n1406), .S1(
        n1410), .Y(n1134) );
  MX4X1 U502 ( .A(\regs[0][4] ), .B(\regs[1][4] ), .C(\regs[2][4] ), .D(
        \regs[3][4] ), .S0(n1440), .S1(n1416), .Y(n1133) );
  MX4X1 U503 ( .A(\regs[8][4] ), .B(\regs[9][4] ), .C(\regs[10][4] ), .D(
        \regs[11][4] ), .S0(n1440), .S1(n1416), .Y(n1131) );
  MX4X1 U504 ( .A(\regs[4][4] ), .B(\regs[5][4] ), .C(\regs[6][4] ), .D(
        \regs[7][4] ), .S0(n1440), .S1(n1416), .Y(n1132) );
  MX4X1 U505 ( .A(n1143), .B(n1141), .C(n1142), .D(n1140), .S0(n1406), .S1(
        n1410), .Y(n1144) );
  MX4X1 U506 ( .A(\regs[0][5] ), .B(\regs[1][5] ), .C(\regs[2][5] ), .D(
        \regs[3][5] ), .S0(n1441), .S1(n1417), .Y(n1143) );
  MX4X1 U507 ( .A(\regs[8][5] ), .B(\regs[9][5] ), .C(\regs[10][5] ), .D(
        \regs[11][5] ), .S0(n1441), .S1(n1417), .Y(n1141) );
  MX4X1 U508 ( .A(\regs[4][5] ), .B(\regs[5][5] ), .C(\regs[6][5] ), .D(
        \regs[7][5] ), .S0(n1441), .S1(n1417), .Y(n1142) );
  MX4X1 U509 ( .A(n1153), .B(n1151), .C(n1152), .D(n1150), .S0(n1406), .S1(
        n1410), .Y(n1154) );
  MX4X1 U510 ( .A(\regs[0][6] ), .B(\regs[1][6] ), .C(\regs[2][6] ), .D(
        \regs[3][6] ), .S0(n1442), .S1(n1418), .Y(n1153) );
  MX4X1 U511 ( .A(\regs[8][6] ), .B(\regs[9][6] ), .C(\regs[10][6] ), .D(
        \regs[11][6] ), .S0(n1442), .S1(n1418), .Y(n1151) );
  MX4X1 U512 ( .A(\regs[4][6] ), .B(\regs[5][6] ), .C(\regs[6][6] ), .D(
        \regs[7][6] ), .S0(n1442), .S1(n1418), .Y(n1152) );
  MX4X1 U513 ( .A(n1163), .B(n1161), .C(n1162), .D(n1160), .S0(n1406), .S1(
        n1410), .Y(n1164) );
  MX4X1 U514 ( .A(\regs[0][7] ), .B(\regs[1][7] ), .C(\regs[2][7] ), .D(
        \regs[3][7] ), .S0(n1442), .S1(n1418), .Y(n1163) );
  MX4X1 U515 ( .A(\regs[8][7] ), .B(\regs[9][7] ), .C(\regs[10][7] ), .D(
        \regs[11][7] ), .S0(n1442), .S1(n1418), .Y(n1161) );
  MX4X1 U516 ( .A(\regs[4][7] ), .B(\regs[5][7] ), .C(\regs[6][7] ), .D(
        \regs[7][7] ), .S0(n1442), .S1(n1418), .Y(n1162) );
  MX4X1 U517 ( .A(n1173), .B(n1171), .C(n1172), .D(n1170), .S0(N15), .S1(n1410), .Y(n1174) );
  MX4X1 U518 ( .A(\regs[0][8] ), .B(\regs[1][8] ), .C(\regs[2][8] ), .D(
        \regs[3][8] ), .S0(n1443), .S1(n1419), .Y(n1173) );
  MX4X1 U519 ( .A(\regs[8][8] ), .B(\regs[9][8] ), .C(\regs[10][8] ), .D(
        \regs[11][8] ), .S0(n1443), .S1(n1419), .Y(n1171) );
  MX4X1 U520 ( .A(\regs[4][8] ), .B(\regs[5][8] ), .C(\regs[6][8] ), .D(
        \regs[7][8] ), .S0(n1443), .S1(n1419), .Y(n1172) );
  MX4X1 U521 ( .A(n1183), .B(n1181), .C(n1182), .D(n1180), .S0(n1406), .S1(
        n1410), .Y(n1184) );
  MX4X1 U522 ( .A(\regs[0][9] ), .B(\regs[1][9] ), .C(\regs[2][9] ), .D(
        \regs[3][9] ), .S0(n1444), .S1(n1420), .Y(n1183) );
  MX4X1 U523 ( .A(\regs[8][9] ), .B(\regs[9][9] ), .C(\regs[10][9] ), .D(
        \regs[11][9] ), .S0(n1444), .S1(n1420), .Y(n1181) );
  MX4X1 U524 ( .A(\regs[4][9] ), .B(\regs[5][9] ), .C(\regs[6][9] ), .D(
        \regs[7][9] ), .S0(n1444), .S1(n1420), .Y(n1182) );
  MX4X1 U525 ( .A(n1193), .B(n1191), .C(n1192), .D(n1190), .S0(N15), .S1(n1410), .Y(n1194) );
  MX4X1 U526 ( .A(\regs[0][10] ), .B(\regs[1][10] ), .C(\regs[2][10] ), .D(
        \regs[3][10] ), .S0(n1444), .S1(n1420), .Y(n1193) );
  MX4X1 U527 ( .A(\regs[8][10] ), .B(\regs[9][10] ), .C(\regs[10][10] ), .D(
        \regs[11][10] ), .S0(n1444), .S1(n1420), .Y(n1191) );
  MX4X1 U528 ( .A(\regs[4][10] ), .B(\regs[5][10] ), .C(\regs[6][10] ), .D(
        \regs[7][10] ), .S0(n1444), .S1(n1420), .Y(n1192) );
  MX4X1 U529 ( .A(n1203), .B(n1201), .C(n1202), .D(n1200), .S0(n1407), .S1(
        n1410), .Y(n1204) );
  MX4X1 U530 ( .A(\regs[0][11] ), .B(\regs[1][11] ), .C(\regs[2][11] ), .D(
        \regs[3][11] ), .S0(n1445), .S1(n1421), .Y(n1203) );
  MX4X1 U531 ( .A(\regs[8][11] ), .B(\regs[9][11] ), .C(\regs[10][11] ), .D(
        \regs[11][11] ), .S0(n1445), .S1(n1421), .Y(n1201) );
  MX4X1 U532 ( .A(\regs[4][11] ), .B(\regs[5][11] ), .C(\regs[6][11] ), .D(
        \regs[7][11] ), .S0(n1445), .S1(n1421), .Y(n1202) );
  MX4X1 U533 ( .A(n1213), .B(n1211), .C(n1212), .D(n1210), .S0(N15), .S1(n1410), .Y(n1214) );
  MX4X1 U534 ( .A(\regs[0][12] ), .B(\regs[1][12] ), .C(\regs[2][12] ), .D(
        \regs[3][12] ), .S0(n1446), .S1(n1422), .Y(n1213) );
  MX4X1 U535 ( .A(\regs[8][12] ), .B(\regs[9][12] ), .C(\regs[10][12] ), .D(
        \regs[11][12] ), .S0(n1446), .S1(n1422), .Y(n1211) );
  MX4X1 U536 ( .A(\regs[4][12] ), .B(\regs[5][12] ), .C(\regs[6][12] ), .D(
        \regs[7][12] ), .S0(n1446), .S1(n1422), .Y(n1212) );
  MX4X1 U537 ( .A(n1223), .B(n1221), .C(n1222), .D(n1220), .S0(n1407), .S1(
        n1410), .Y(n1224) );
  MX4X1 U538 ( .A(\regs[0][13] ), .B(\regs[1][13] ), .C(\regs[2][13] ), .D(
        \regs[3][13] ), .S0(n1446), .S1(n1422), .Y(n1223) );
  MX4X1 U539 ( .A(\regs[8][13] ), .B(\regs[9][13] ), .C(\regs[10][13] ), .D(
        \regs[11][13] ), .S0(n1446), .S1(n1422), .Y(n1221) );
  MX4X1 U540 ( .A(\regs[4][13] ), .B(\regs[5][13] ), .C(\regs[6][13] ), .D(
        \regs[7][13] ), .S0(n1446), .S1(n1422), .Y(n1222) );
  MX4X1 U541 ( .A(n1233), .B(n1231), .C(n1232), .D(n1230), .S0(n1407), .S1(N14), .Y(n1234) );
  MX4X1 U542 ( .A(\regs[0][14] ), .B(\regs[1][14] ), .C(\regs[2][14] ), .D(
        \regs[3][14] ), .S0(n1447), .S1(n1423), .Y(n1233) );
  MX4X1 U543 ( .A(\regs[8][14] ), .B(\regs[9][14] ), .C(\regs[10][14] ), .D(
        \regs[11][14] ), .S0(n1447), .S1(n1423), .Y(n1231) );
  MX4X1 U544 ( .A(\regs[4][14] ), .B(\regs[5][14] ), .C(\regs[6][14] ), .D(
        \regs[7][14] ), .S0(n1447), .S1(n1423), .Y(n1232) );
  MX4X1 U545 ( .A(n1243), .B(n1241), .C(n1242), .D(n1240), .S0(n1407), .S1(N14), .Y(n1244) );
  MX4X1 U546 ( .A(\regs[0][15] ), .B(\regs[1][15] ), .C(\regs[2][15] ), .D(
        \regs[3][15] ), .S0(n1448), .S1(n1424), .Y(n1243) );
  MX4X1 U547 ( .A(\regs[8][15] ), .B(\regs[9][15] ), .C(\regs[10][15] ), .D(
        \regs[11][15] ), .S0(n1448), .S1(n1424), .Y(n1241) );
  MX4X1 U548 ( .A(\regs[4][15] ), .B(\regs[5][15] ), .C(\regs[6][15] ), .D(
        \regs[7][15] ), .S0(n1448), .S1(n1424), .Y(n1242) );
  MX4X1 U549 ( .A(n1253), .B(n1251), .C(n1252), .D(n1250), .S0(n1407), .S1(N14), .Y(n1254) );
  MX4X1 U550 ( .A(\regs[0][16] ), .B(\regs[1][16] ), .C(\regs[2][16] ), .D(
        \regs[3][16] ), .S0(n1448), .S1(n1424), .Y(n1253) );
  MX4X1 U551 ( .A(\regs[8][16] ), .B(\regs[9][16] ), .C(\regs[10][16] ), .D(
        \regs[11][16] ), .S0(n1448), .S1(n1424), .Y(n1251) );
  MX4X1 U552 ( .A(\regs[4][16] ), .B(\regs[5][16] ), .C(\regs[6][16] ), .D(
        \regs[7][16] ), .S0(n1448), .S1(n1424), .Y(n1252) );
  MX4X1 U553 ( .A(n1263), .B(n1261), .C(n1262), .D(n1260), .S0(n1407), .S1(
        n1410), .Y(n1264) );
  MX4X1 U554 ( .A(\regs[0][17] ), .B(\regs[1][17] ), .C(\regs[2][17] ), .D(
        \regs[3][17] ), .S0(n1449), .S1(n1425), .Y(n1263) );
  MX4X1 U555 ( .A(\regs[8][17] ), .B(\regs[9][17] ), .C(\regs[10][17] ), .D(
        \regs[11][17] ), .S0(n1449), .S1(n1425), .Y(n1261) );
  MX4X1 U556 ( .A(\regs[4][17] ), .B(\regs[5][17] ), .C(\regs[6][17] ), .D(
        \regs[7][17] ), .S0(n1449), .S1(n1425), .Y(n1262) );
  MX4X1 U557 ( .A(n1273), .B(n1271), .C(n1272), .D(n1270), .S0(n1407), .S1(N14), .Y(n1274) );
  MX4X1 U558 ( .A(\regs[0][18] ), .B(\regs[1][18] ), .C(\regs[2][18] ), .D(
        \regs[3][18] ), .S0(n1450), .S1(n1426), .Y(n1273) );
  MX4X1 U559 ( .A(\regs[8][18] ), .B(\regs[9][18] ), .C(\regs[10][18] ), .D(
        \regs[11][18] ), .S0(n1450), .S1(n1426), .Y(n1271) );
  MX4X1 U560 ( .A(\regs[4][18] ), .B(\regs[5][18] ), .C(\regs[6][18] ), .D(
        \regs[7][18] ), .S0(n1450), .S1(n1426), .Y(n1272) );
  MX4X1 U561 ( .A(n1283), .B(n1281), .C(n1282), .D(n1280), .S0(n1407), .S1(N14), .Y(n1284) );
  MX4X1 U562 ( .A(\regs[0][19] ), .B(\regs[1][19] ), .C(\regs[2][19] ), .D(
        \regs[3][19] ), .S0(n1450), .S1(n1426), .Y(n1283) );
  MX4X1 U563 ( .A(\regs[8][19] ), .B(\regs[9][19] ), .C(\regs[10][19] ), .D(
        \regs[11][19] ), .S0(n1450), .S1(n1426), .Y(n1281) );
  MX4X1 U564 ( .A(\regs[4][19] ), .B(\regs[5][19] ), .C(\regs[6][19] ), .D(
        \regs[7][19] ), .S0(n1450), .S1(n1426), .Y(n1282) );
  MX4X1 U565 ( .A(n1293), .B(n1291), .C(n1292), .D(n1290), .S0(n1408), .S1(N14), .Y(n1294) );
  MX4X1 U566 ( .A(\regs[0][20] ), .B(\regs[1][20] ), .C(\regs[2][20] ), .D(
        \regs[3][20] ), .S0(n1451), .S1(n1427), .Y(n1293) );
  MX4X1 U567 ( .A(\regs[8][20] ), .B(\regs[9][20] ), .C(\regs[10][20] ), .D(
        \regs[11][20] ), .S0(n1451), .S1(n1427), .Y(n1291) );
  MX4X1 U568 ( .A(\regs[4][20] ), .B(\regs[5][20] ), .C(\regs[6][20] ), .D(
        \regs[7][20] ), .S0(n1451), .S1(n1427), .Y(n1292) );
  MX4X1 U569 ( .A(n1303), .B(n1301), .C(n1302), .D(n1300), .S0(N15), .S1(N14), 
        .Y(n1304) );
  MX4X1 U570 ( .A(\regs[0][21] ), .B(\regs[1][21] ), .C(\regs[2][21] ), .D(
        \regs[3][21] ), .S0(n1452), .S1(n1428), .Y(n1303) );
  MX4X1 U571 ( .A(\regs[8][21] ), .B(\regs[9][21] ), .C(\regs[10][21] ), .D(
        \regs[11][21] ), .S0(n1452), .S1(n1428), .Y(n1301) );
  MX4X1 U572 ( .A(\regs[4][21] ), .B(\regs[5][21] ), .C(\regs[6][21] ), .D(
        \regs[7][21] ), .S0(n1452), .S1(n1428), .Y(n1302) );
  MX4X1 U573 ( .A(n1313), .B(n1311), .C(n1312), .D(n1310), .S0(N15), .S1(N14), 
        .Y(n1314) );
  MX4X1 U574 ( .A(\regs[0][22] ), .B(\regs[1][22] ), .C(\regs[2][22] ), .D(
        \regs[3][22] ), .S0(n1452), .S1(n1428), .Y(n1313) );
  MX4X1 U575 ( .A(\regs[8][22] ), .B(\regs[9][22] ), .C(\regs[10][22] ), .D(
        \regs[11][22] ), .S0(n1452), .S1(n1428), .Y(n1311) );
  MX4X1 U576 ( .A(\regs[4][22] ), .B(\regs[5][22] ), .C(\regs[6][22] ), .D(
        \regs[7][22] ), .S0(n1452), .S1(n1428), .Y(n1312) );
  MX4X1 U577 ( .A(n1323), .B(n1321), .C(n1322), .D(n1320), .S0(N15), .S1(n1410), .Y(n1324) );
  MX4X1 U578 ( .A(\regs[0][23] ), .B(\regs[1][23] ), .C(\regs[2][23] ), .D(
        \regs[3][23] ), .S0(n1453), .S1(n1429), .Y(n1323) );
  MX4X1 U579 ( .A(\regs[8][23] ), .B(\regs[9][23] ), .C(\regs[10][23] ), .D(
        \regs[11][23] ), .S0(n1453), .S1(n1429), .Y(n1321) );
  MX4X1 U580 ( .A(\regs[4][23] ), .B(\regs[5][23] ), .C(\regs[6][23] ), .D(
        \regs[7][23] ), .S0(n1453), .S1(n1429), .Y(n1322) );
  MX4X1 U581 ( .A(n1333), .B(n1331), .C(n1332), .D(n1330), .S0(n1406), .S1(N14), .Y(n1334) );
  MX4X1 U582 ( .A(\regs[0][24] ), .B(\regs[1][24] ), .C(\regs[2][24] ), .D(
        \regs[3][24] ), .S0(n1454), .S1(n1430), .Y(n1333) );
  MX4X1 U583 ( .A(\regs[8][24] ), .B(\regs[9][24] ), .C(\regs[10][24] ), .D(
        \regs[11][24] ), .S0(n1454), .S1(n1430), .Y(n1331) );
  MX4X1 U584 ( .A(\regs[4][24] ), .B(\regs[5][24] ), .C(\regs[6][24] ), .D(
        \regs[7][24] ), .S0(n1454), .S1(n1430), .Y(n1332) );
  MX4X1 U585 ( .A(n1343), .B(n1341), .C(n1342), .D(n1340), .S0(N15), .S1(n1410), .Y(n1344) );
  MX4X1 U586 ( .A(\regs[0][25] ), .B(\regs[1][25] ), .C(\regs[2][25] ), .D(
        \regs[3][25] ), .S0(n1454), .S1(n1430), .Y(n1343) );
  MX4X1 U587 ( .A(\regs[8][25] ), .B(\regs[9][25] ), .C(\regs[10][25] ), .D(
        \regs[11][25] ), .S0(n1454), .S1(n1430), .Y(n1341) );
  MX4X1 U588 ( .A(\regs[4][25] ), .B(\regs[5][25] ), .C(\regs[6][25] ), .D(
        \regs[7][25] ), .S0(n1454), .S1(n1430), .Y(n1342) );
  MX4X1 U589 ( .A(n1393), .B(n1391), .C(n1392), .D(n1390), .S0(n1408), .S1(N14), .Y(n1394) );
  MX4X1 U590 ( .A(\regs[0][30] ), .B(\regs[1][30] ), .C(\regs[2][30] ), .D(
        \regs[3][30] ), .S0(n1458), .S1(n1434), .Y(n1393) );
  MX4X1 U591 ( .A(\regs[8][30] ), .B(\regs[9][30] ), .C(\regs[10][30] ), .D(
        \regs[11][30] ), .S0(n1458), .S1(n1434), .Y(n1391) );
  MX4X1 U592 ( .A(\regs[4][30] ), .B(\regs[5][30] ), .C(\regs[6][30] ), .D(
        \regs[7][30] ), .S0(n1458), .S1(n1434), .Y(n1392) );
  MX4X1 U593 ( .A(n1403), .B(n1401), .C(n1402), .D(n1400), .S0(n1408), .S1(N14), .Y(n1404) );
  MX4X1 U594 ( .A(\regs[0][31] ), .B(\regs[1][31] ), .C(\regs[2][31] ), .D(
        \regs[3][31] ), .S0(n1458), .S1(n1434), .Y(n1403) );
  MX4X1 U595 ( .A(\regs[8][31] ), .B(\regs[9][31] ), .C(\regs[10][31] ), .D(
        \regs[11][31] ), .S0(n1458), .S1(n1434), .Y(n1401) );
  MX4X1 U596 ( .A(\regs[4][31] ), .B(\regs[5][31] ), .C(\regs[6][31] ), .D(
        \regs[7][31] ), .S0(n1458), .S1(n1434), .Y(n1402) );
  MX4X1 U597 ( .A(\regs[20][26] ), .B(\regs[21][26] ), .C(\regs[22][26] ), .D(
        \regs[23][26] ), .S0(n1455), .S1(n1431), .Y(n1347) );
  MX4X1 U598 ( .A(\regs[4][26] ), .B(\regs[5][26] ), .C(\regs[6][26] ), .D(
        \regs[7][26] ), .S0(n1455), .S1(n1431), .Y(n1352) );
  MX4X1 U599 ( .A(\regs[20][27] ), .B(\regs[21][27] ), .C(\regs[22][27] ), .D(
        \regs[23][27] ), .S0(n1455), .S1(n1431), .Y(n1357) );
  MX4X1 U600 ( .A(\regs[4][27] ), .B(\regs[5][27] ), .C(\regs[6][27] ), .D(
        \regs[7][27] ), .S0(n1456), .S1(n1432), .Y(n1362) );
  MX4X1 U601 ( .A(\regs[20][28] ), .B(\regs[21][28] ), .C(\regs[22][28] ), .D(
        \regs[23][28] ), .S0(n1456), .S1(n1432), .Y(n1367) );
  MX4X1 U602 ( .A(\regs[4][28] ), .B(\regs[5][28] ), .C(\regs[6][28] ), .D(
        \regs[7][28] ), .S0(n1456), .S1(n1432), .Y(n1372) );
  MX4X1 U603 ( .A(\regs[20][29] ), .B(\regs[21][29] ), .C(\regs[22][29] ), .D(
        \regs[23][29] ), .S0(n1457), .S1(n1433), .Y(n1377) );
  MX4X1 U604 ( .A(\regs[4][29] ), .B(\regs[5][29] ), .C(\regs[6][29] ), .D(
        \regs[7][29] ), .S0(n1457), .S1(n1433), .Y(n1382) );
  MX4X1 U605 ( .A(\regs[16][26] ), .B(\regs[17][26] ), .C(\regs[18][26] ), .D(
        \regs[19][26] ), .S0(n1455), .S1(n1431), .Y(n1348) );
  MX4X1 U606 ( .A(\regs[16][27] ), .B(\regs[17][27] ), .C(\regs[18][27] ), .D(
        \regs[19][27] ), .S0(n1455), .S1(n1431), .Y(n1358) );
  MX4X1 U607 ( .A(\regs[16][28] ), .B(\regs[17][28] ), .C(\regs[18][28] ), .D(
        \regs[19][28] ), .S0(n1456), .S1(n1432), .Y(n1368) );
  MX4X1 U608 ( .A(\regs[16][29] ), .B(\regs[17][29] ), .C(\regs[18][29] ), .D(
        \regs[19][29] ), .S0(n1457), .S1(n1433), .Y(n1378) );
  MX4X1 U609 ( .A(\regs[12][0] ), .B(\regs[13][0] ), .C(\regs[14][0] ), .D(
        \regs[15][0] ), .S0(n2183), .S1(n2158), .Y(n1835) );
  MX4X1 U610 ( .A(\regs[28][0] ), .B(\regs[29][0] ), .C(\regs[30][0] ), .D(
        \regs[31][0] ), .S0(n2188), .S1(n2174), .Y(n1830) );
  MX4X1 U611 ( .A(\regs[28][1] ), .B(\regs[29][1] ), .C(\regs[30][1] ), .D(
        \regs[31][1] ), .S0(n2183), .S1(n2158), .Y(n1840) );
  MX4X1 U612 ( .A(\regs[12][1] ), .B(\regs[13][1] ), .C(\regs[14][1] ), .D(
        \regs[15][1] ), .S0(n2183), .S1(n2158), .Y(n1845) );
  MX4X1 U613 ( .A(\regs[28][2] ), .B(\regs[29][2] ), .C(\regs[30][2] ), .D(
        \regs[31][2] ), .S0(n2184), .S1(n2159), .Y(n1850) );
  MX4X1 U614 ( .A(\regs[12][2] ), .B(\regs[13][2] ), .C(\regs[14][2] ), .D(
        \regs[15][2] ), .S0(n2184), .S1(n2159), .Y(n1855) );
  MX4X1 U615 ( .A(\regs[28][3] ), .B(\regs[29][3] ), .C(\regs[30][3] ), .D(
        \regs[31][3] ), .S0(n2184), .S1(n2159), .Y(n1860) );
  MX4X1 U616 ( .A(\regs[12][3] ), .B(\regs[13][3] ), .C(\regs[14][3] ), .D(
        \regs[15][3] ), .S0(n2185), .S1(n2160), .Y(n1865) );
  MX4X1 U617 ( .A(\regs[28][4] ), .B(\regs[29][4] ), .C(\regs[30][4] ), .D(
        \regs[31][4] ), .S0(n2185), .S1(n2160), .Y(n1870) );
  MX4X1 U618 ( .A(\regs[12][4] ), .B(\regs[13][4] ), .C(\regs[14][4] ), .D(
        \regs[15][4] ), .S0(n2185), .S1(n2160), .Y(n1875) );
  MX4X1 U619 ( .A(\regs[28][5] ), .B(\regs[29][5] ), .C(\regs[30][5] ), .D(
        \regs[31][5] ), .S0(n2186), .S1(n2161), .Y(n1880) );
  MX4X1 U620 ( .A(\regs[12][5] ), .B(\regs[13][5] ), .C(\regs[14][5] ), .D(
        \regs[15][5] ), .S0(n2186), .S1(n2161), .Y(n1885) );
  MX4X1 U621 ( .A(\regs[28][6] ), .B(\regs[29][6] ), .C(\regs[30][6] ), .D(
        \regs[31][6] ), .S0(n2186), .S1(n2161), .Y(n1890) );
  MX4X1 U622 ( .A(\regs[12][6] ), .B(\regs[13][6] ), .C(\regs[14][6] ), .D(
        \regs[15][6] ), .S0(n2187), .S1(n2162), .Y(n1895) );
  MX4X1 U623 ( .A(\regs[28][7] ), .B(\regs[29][7] ), .C(\regs[30][7] ), .D(
        \regs[31][7] ), .S0(n2187), .S1(n2162), .Y(n1900) );
  MX4X1 U624 ( .A(\regs[12][7] ), .B(\regs[13][7] ), .C(\regs[14][7] ), .D(
        \regs[15][7] ), .S0(n2187), .S1(n2162), .Y(n1905) );
  MX4X1 U625 ( .A(\regs[28][8] ), .B(\regs[29][8] ), .C(\regs[30][8] ), .D(
        \regs[31][8] ), .S0(n2188), .S1(n2163), .Y(n1910) );
  MX4X1 U626 ( .A(\regs[12][8] ), .B(\regs[13][8] ), .C(\regs[14][8] ), .D(
        \regs[15][8] ), .S0(n2188), .S1(n2163), .Y(n1915) );
  MX4X1 U627 ( .A(\regs[28][9] ), .B(\regs[29][9] ), .C(\regs[30][9] ), .D(
        \regs[31][9] ), .S0(n2188), .S1(n2163), .Y(n1920) );
  MX4X1 U628 ( .A(\regs[12][9] ), .B(\regs[13][9] ), .C(\regs[14][9] ), .D(
        \regs[15][9] ), .S0(n2189), .S1(n2164), .Y(n1925) );
  MX4X1 U629 ( .A(\regs[28][10] ), .B(\regs[29][10] ), .C(\regs[30][10] ), .D(
        \regs[31][10] ), .S0(n2189), .S1(n2164), .Y(n1930) );
  MX4X1 U630 ( .A(\regs[12][10] ), .B(\regs[13][10] ), .C(\regs[14][10] ), .D(
        \regs[15][10] ), .S0(n2189), .S1(n2164), .Y(n1935) );
  MX4X1 U631 ( .A(\regs[28][11] ), .B(\regs[29][11] ), .C(\regs[30][11] ), .D(
        \regs[31][11] ), .S0(n2190), .S1(n2165), .Y(n1940) );
  MX4X1 U632 ( .A(\regs[12][11] ), .B(\regs[13][11] ), .C(\regs[14][11] ), .D(
        \regs[15][11] ), .S0(n2190), .S1(n2165), .Y(n1945) );
  MX4X1 U633 ( .A(\regs[28][12] ), .B(\regs[29][12] ), .C(\regs[30][12] ), .D(
        \regs[31][12] ), .S0(n2190), .S1(n2165), .Y(n1950) );
  MX4X1 U634 ( .A(\regs[12][12] ), .B(\regs[13][12] ), .C(\regs[14][12] ), .D(
        \regs[15][12] ), .S0(n2191), .S1(n2166), .Y(n1955) );
  MX4X1 U635 ( .A(\regs[28][13] ), .B(\regs[29][13] ), .C(\regs[30][13] ), .D(
        \regs[31][13] ), .S0(n2191), .S1(n2166), .Y(n1960) );
  MX4X1 U636 ( .A(\regs[12][13] ), .B(\regs[13][13] ), .C(\regs[14][13] ), .D(
        \regs[15][13] ), .S0(n2191), .S1(n2166), .Y(n1965) );
  MX4X1 U637 ( .A(\regs[28][14] ), .B(\regs[29][14] ), .C(\regs[30][14] ), .D(
        \regs[31][14] ), .S0(n2192), .S1(n2167), .Y(n1970) );
  MX4X1 U638 ( .A(\regs[12][14] ), .B(\regs[13][14] ), .C(\regs[14][14] ), .D(
        \regs[15][14] ), .S0(n2192), .S1(n2167), .Y(n1975) );
  MX4X1 U639 ( .A(\regs[28][15] ), .B(\regs[29][15] ), .C(\regs[30][15] ), .D(
        \regs[31][15] ), .S0(n2192), .S1(n2167), .Y(n1980) );
  MX4X1 U640 ( .A(\regs[12][15] ), .B(\regs[13][15] ), .C(\regs[14][15] ), .D(
        \regs[15][15] ), .S0(n2193), .S1(n2168), .Y(n1985) );
  MX4X1 U641 ( .A(\regs[28][16] ), .B(\regs[29][16] ), .C(\regs[30][16] ), .D(
        \regs[31][16] ), .S0(n2193), .S1(n2168), .Y(n1990) );
  MX4X1 U642 ( .A(\regs[12][16] ), .B(\regs[13][16] ), .C(\regs[14][16] ), .D(
        \regs[15][16] ), .S0(n2193), .S1(n2168), .Y(n1995) );
  MX4X1 U643 ( .A(\regs[28][17] ), .B(\regs[29][17] ), .C(\regs[30][17] ), .D(
        \regs[31][17] ), .S0(n2194), .S1(n2169), .Y(n2000) );
  MX4X1 U644 ( .A(\regs[12][17] ), .B(\regs[13][17] ), .C(\regs[14][17] ), .D(
        \regs[15][17] ), .S0(n2194), .S1(n2169), .Y(n2005) );
  MX4X1 U645 ( .A(\regs[28][18] ), .B(\regs[29][18] ), .C(\regs[30][18] ), .D(
        \regs[31][18] ), .S0(n2194), .S1(n2169), .Y(n2010) );
  MX4X1 U646 ( .A(\regs[12][18] ), .B(\regs[13][18] ), .C(\regs[14][18] ), .D(
        \regs[15][18] ), .S0(n2195), .S1(n2170), .Y(n2015) );
  MX4X1 U647 ( .A(\regs[28][19] ), .B(\regs[29][19] ), .C(\regs[30][19] ), .D(
        \regs[31][19] ), .S0(n2195), .S1(n2170), .Y(n2020) );
  MX4X1 U648 ( .A(\regs[12][19] ), .B(\regs[13][19] ), .C(\regs[14][19] ), .D(
        \regs[15][19] ), .S0(n2195), .S1(n2170), .Y(n2025) );
  MX4X1 U649 ( .A(\regs[28][20] ), .B(\regs[29][20] ), .C(\regs[30][20] ), .D(
        \regs[31][20] ), .S0(n2196), .S1(n2171), .Y(n2030) );
  MX4X1 U650 ( .A(\regs[12][20] ), .B(\regs[13][20] ), .C(\regs[14][20] ), .D(
        \regs[15][20] ), .S0(n2196), .S1(n2171), .Y(n2035) );
  MX4X1 U651 ( .A(\regs[28][21] ), .B(\regs[29][21] ), .C(\regs[30][21] ), .D(
        \regs[31][21] ), .S0(n2196), .S1(n2171), .Y(n2040) );
  MX4X1 U652 ( .A(\regs[12][21] ), .B(\regs[13][21] ), .C(\regs[14][21] ), .D(
        \regs[15][21] ), .S0(n2197), .S1(n2172), .Y(n2045) );
  MX4X1 U653 ( .A(\regs[28][22] ), .B(\regs[29][22] ), .C(\regs[30][22] ), .D(
        \regs[31][22] ), .S0(n2197), .S1(n2172), .Y(n2050) );
  MX4X1 U654 ( .A(\regs[12][22] ), .B(\regs[13][22] ), .C(\regs[14][22] ), .D(
        \regs[15][22] ), .S0(n2197), .S1(n2172), .Y(n2055) );
  MX4X1 U655 ( .A(\regs[28][23] ), .B(\regs[29][23] ), .C(\regs[30][23] ), .D(
        \regs[31][23] ), .S0(n2198), .S1(n2173), .Y(n2060) );
  MX4X1 U656 ( .A(\regs[12][23] ), .B(\regs[13][23] ), .C(\regs[14][23] ), .D(
        \regs[15][23] ), .S0(n2198), .S1(n2173), .Y(n2065) );
  MX4X1 U657 ( .A(\regs[28][24] ), .B(\regs[29][24] ), .C(\regs[30][24] ), .D(
        \regs[31][24] ), .S0(n2198), .S1(n2173), .Y(n2070) );
  MX4X1 U658 ( .A(\regs[12][24] ), .B(\regs[13][24] ), .C(\regs[14][24] ), .D(
        \regs[15][24] ), .S0(n2199), .S1(n2174), .Y(n2075) );
  MX4X1 U659 ( .A(\regs[28][25] ), .B(\regs[29][25] ), .C(\regs[30][25] ), .D(
        \regs[31][25] ), .S0(n2199), .S1(n2174), .Y(n2080) );
  MX4X1 U660 ( .A(\regs[12][25] ), .B(\regs[13][25] ), .C(\regs[14][25] ), .D(
        \regs[15][25] ), .S0(n2199), .S1(n2174), .Y(n2085) );
  MX4X1 U661 ( .A(\regs[28][26] ), .B(\regs[29][26] ), .C(\regs[30][26] ), .D(
        \regs[31][26] ), .S0(n2200), .S1(n2175), .Y(n2090) );
  MX4X1 U662 ( .A(\regs[12][26] ), .B(\regs[13][26] ), .C(\regs[14][26] ), .D(
        \regs[15][26] ), .S0(n2200), .S1(n2175), .Y(n2095) );
  MX4X1 U663 ( .A(\regs[28][27] ), .B(\regs[29][27] ), .C(\regs[30][27] ), .D(
        \regs[31][27] ), .S0(n2200), .S1(n2175), .Y(n2100) );
  MX4X1 U664 ( .A(\regs[12][27] ), .B(\regs[13][27] ), .C(\regs[14][27] ), .D(
        \regs[15][27] ), .S0(n2201), .S1(n2176), .Y(n2105) );
  MX4X1 U665 ( .A(\regs[28][28] ), .B(\regs[29][28] ), .C(\regs[30][28] ), .D(
        \regs[31][28] ), .S0(n2201), .S1(n2176), .Y(n2110) );
  MX4X1 U666 ( .A(\regs[12][28] ), .B(\regs[13][28] ), .C(\regs[14][28] ), .D(
        \regs[15][28] ), .S0(n2201), .S1(n2176), .Y(n2115) );
  MX4X1 U667 ( .A(\regs[28][29] ), .B(\regs[29][29] ), .C(\regs[30][29] ), .D(
        \regs[31][29] ), .S0(n2202), .S1(n2177), .Y(n2120) );
  MX4X1 U668 ( .A(\regs[12][29] ), .B(\regs[13][29] ), .C(\regs[14][29] ), .D(
        \regs[15][29] ), .S0(n2202), .S1(n2177), .Y(n2125) );
  MX4X1 U669 ( .A(\regs[28][30] ), .B(\regs[29][30] ), .C(\regs[30][30] ), .D(
        \regs[31][30] ), .S0(n2202), .S1(n2177), .Y(n2130) );
  MX4X1 U670 ( .A(\regs[12][30] ), .B(\regs[13][30] ), .C(\regs[14][30] ), .D(
        \regs[15][30] ), .S0(n2203), .S1(n2178), .Y(n2135) );
  MX4X1 U671 ( .A(\regs[28][31] ), .B(\regs[29][31] ), .C(\regs[30][31] ), .D(
        \regs[31][31] ), .S0(n2203), .S1(n2178), .Y(n2140) );
  MX4X1 U672 ( .A(\regs[12][31] ), .B(\regs[13][31] ), .C(\regs[14][31] ), .D(
        \regs[15][31] ), .S0(n2203), .S1(n2178), .Y(n2145) );
  MX4X1 U673 ( .A(\regs[12][0] ), .B(\regs[13][0] ), .C(\regs[14][0] ), .D(
        \regs[15][0] ), .S0(n1438), .S1(n1414), .Y(n53) );
  MX4X1 U674 ( .A(\regs[28][0] ), .B(\regs[29][0] ), .C(\regs[30][0] ), .D(
        \regs[31][0] ), .S0(n1443), .S1(n1421), .Y(n45) );
  MX4X1 U675 ( .A(\regs[28][1] ), .B(\regs[29][1] ), .C(\regs[30][1] ), .D(
        \regs[31][1] ), .S0(n1438), .S1(n1414), .Y(n60) );
  MX4X1 U676 ( .A(\regs[12][1] ), .B(\regs[13][1] ), .C(\regs[14][1] ), .D(
        \regs[15][1] ), .S0(n1438), .S1(n1414), .Y(n72) );
  MX4X1 U677 ( .A(\regs[28][2] ), .B(\regs[29][2] ), .C(\regs[30][2] ), .D(
        \regs[31][2] ), .S0(n1439), .S1(n1415), .Y(n79) );
  MX4X1 U678 ( .A(\regs[12][2] ), .B(\regs[13][2] ), .C(\regs[14][2] ), .D(
        \regs[15][2] ), .S0(n1439), .S1(n1415), .Y(n1110) );
  MX4X1 U679 ( .A(\regs[28][3] ), .B(\regs[29][3] ), .C(\regs[30][3] ), .D(
        \regs[31][3] ), .S0(n1439), .S1(n1415), .Y(n1115) );
  MX4X1 U680 ( .A(\regs[12][3] ), .B(\regs[13][3] ), .C(\regs[14][3] ), .D(
        \regs[15][3] ), .S0(n1440), .S1(n1416), .Y(n1120) );
  MX4X1 U681 ( .A(\regs[28][4] ), .B(\regs[29][4] ), .C(\regs[30][4] ), .D(
        \regs[31][4] ), .S0(n1440), .S1(n1416), .Y(n1125) );
  MX4X1 U682 ( .A(\regs[12][4] ), .B(\regs[13][4] ), .C(\regs[14][4] ), .D(
        \regs[15][4] ), .S0(n1440), .S1(n1416), .Y(n1130) );
  MX4X1 U683 ( .A(\regs[28][5] ), .B(\regs[29][5] ), .C(\regs[30][5] ), .D(
        \regs[31][5] ), .S0(n1441), .S1(n1417), .Y(n1135) );
  MX4X1 U684 ( .A(\regs[12][5] ), .B(\regs[13][5] ), .C(\regs[14][5] ), .D(
        \regs[15][5] ), .S0(n1441), .S1(n1417), .Y(n1140) );
  MX4X1 U685 ( .A(\regs[28][6] ), .B(\regs[29][6] ), .C(\regs[30][6] ), .D(
        \regs[31][6] ), .S0(n1441), .S1(n1417), .Y(n1145) );
  MX4X1 U686 ( .A(\regs[12][6] ), .B(\regs[13][6] ), .C(\regs[14][6] ), .D(
        \regs[15][6] ), .S0(n1442), .S1(n1418), .Y(n1150) );
  MX4X1 U687 ( .A(\regs[28][7] ), .B(\regs[29][7] ), .C(\regs[30][7] ), .D(
        \regs[31][7] ), .S0(n1442), .S1(n1418), .Y(n1155) );
  MX4X1 U688 ( .A(\regs[12][7] ), .B(\regs[13][7] ), .C(\regs[14][7] ), .D(
        \regs[15][7] ), .S0(n1442), .S1(n1418), .Y(n1160) );
  MX4X1 U689 ( .A(\regs[28][8] ), .B(\regs[29][8] ), .C(\regs[30][8] ), .D(
        \regs[31][8] ), .S0(n1443), .S1(n1419), .Y(n1165) );
  MX4X1 U690 ( .A(\regs[12][8] ), .B(\regs[13][8] ), .C(\regs[14][8] ), .D(
        \regs[15][8] ), .S0(n1443), .S1(n1419), .Y(n1170) );
  MX4X1 U691 ( .A(\regs[28][9] ), .B(\regs[29][9] ), .C(\regs[30][9] ), .D(
        \regs[31][9] ), .S0(n1443), .S1(n1419), .Y(n1175) );
  MX4X1 U692 ( .A(\regs[12][9] ), .B(\regs[13][9] ), .C(\regs[14][9] ), .D(
        \regs[15][9] ), .S0(n1444), .S1(n1420), .Y(n1180) );
  MX4X1 U693 ( .A(\regs[28][10] ), .B(\regs[29][10] ), .C(\regs[30][10] ), .D(
        \regs[31][10] ), .S0(n1444), .S1(n1420), .Y(n1185) );
  MX4X1 U694 ( .A(\regs[12][10] ), .B(\regs[13][10] ), .C(\regs[14][10] ), .D(
        \regs[15][10] ), .S0(n1444), .S1(n1420), .Y(n1190) );
  MX4X1 U695 ( .A(\regs[28][11] ), .B(\regs[29][11] ), .C(\regs[30][11] ), .D(
        \regs[31][11] ), .S0(n1445), .S1(n1421), .Y(n1195) );
  MX4X1 U696 ( .A(\regs[12][11] ), .B(\regs[13][11] ), .C(\regs[14][11] ), .D(
        \regs[15][11] ), .S0(n1445), .S1(n1421), .Y(n1200) );
  MX4X1 U697 ( .A(\regs[28][12] ), .B(\regs[29][12] ), .C(\regs[30][12] ), .D(
        \regs[31][12] ), .S0(n1445), .S1(n1421), .Y(n1205) );
  MX4X1 U698 ( .A(\regs[12][12] ), .B(\regs[13][12] ), .C(\regs[14][12] ), .D(
        \regs[15][12] ), .S0(n1446), .S1(n1422), .Y(n1210) );
  MX4X1 U699 ( .A(\regs[28][13] ), .B(\regs[29][13] ), .C(\regs[30][13] ), .D(
        \regs[31][13] ), .S0(n1446), .S1(n1422), .Y(n1215) );
  MX4X1 U700 ( .A(\regs[12][13] ), .B(\regs[13][13] ), .C(\regs[14][13] ), .D(
        \regs[15][13] ), .S0(n1446), .S1(n1422), .Y(n1220) );
  MX4X1 U701 ( .A(\regs[28][14] ), .B(\regs[29][14] ), .C(\regs[30][14] ), .D(
        \regs[31][14] ), .S0(n1447), .S1(n1423), .Y(n1225) );
  MX4X1 U702 ( .A(\regs[12][14] ), .B(\regs[13][14] ), .C(\regs[14][14] ), .D(
        \regs[15][14] ), .S0(n1447), .S1(n1423), .Y(n1230) );
  MX4X1 U703 ( .A(\regs[28][15] ), .B(\regs[29][15] ), .C(\regs[30][15] ), .D(
        \regs[31][15] ), .S0(n1447), .S1(n1423), .Y(n1235) );
  MX4X1 U704 ( .A(\regs[12][15] ), .B(\regs[13][15] ), .C(\regs[14][15] ), .D(
        \regs[15][15] ), .S0(n1448), .S1(n1424), .Y(n1240) );
  MX4X1 U705 ( .A(\regs[28][16] ), .B(\regs[29][16] ), .C(\regs[30][16] ), .D(
        \regs[31][16] ), .S0(n1448), .S1(n1424), .Y(n1245) );
  MX4X1 U706 ( .A(\regs[12][16] ), .B(\regs[13][16] ), .C(\regs[14][16] ), .D(
        \regs[15][16] ), .S0(n1448), .S1(n1424), .Y(n1250) );
  MX4X1 U707 ( .A(\regs[28][17] ), .B(\regs[29][17] ), .C(\regs[30][17] ), .D(
        \regs[31][17] ), .S0(n1449), .S1(n1425), .Y(n1255) );
  MX4X1 U708 ( .A(\regs[12][17] ), .B(\regs[13][17] ), .C(\regs[14][17] ), .D(
        \regs[15][17] ), .S0(n1449), .S1(n1425), .Y(n1260) );
  MX4X1 U709 ( .A(\regs[28][18] ), .B(\regs[29][18] ), .C(\regs[30][18] ), .D(
        \regs[31][18] ), .S0(n1449), .S1(n1425), .Y(n1265) );
  MX4X1 U710 ( .A(\regs[12][18] ), .B(\regs[13][18] ), .C(\regs[14][18] ), .D(
        \regs[15][18] ), .S0(n1450), .S1(n1426), .Y(n1270) );
  MX4X1 U711 ( .A(\regs[28][19] ), .B(\regs[29][19] ), .C(\regs[30][19] ), .D(
        \regs[31][19] ), .S0(n1450), .S1(n1426), .Y(n1275) );
  MX4X1 U712 ( .A(\regs[12][19] ), .B(\regs[13][19] ), .C(\regs[14][19] ), .D(
        \regs[15][19] ), .S0(n1450), .S1(n1426), .Y(n1280) );
  MX4X1 U713 ( .A(\regs[28][20] ), .B(\regs[29][20] ), .C(\regs[30][20] ), .D(
        \regs[31][20] ), .S0(n1451), .S1(n1427), .Y(n1285) );
  MX4X1 U714 ( .A(\regs[12][20] ), .B(\regs[13][20] ), .C(\regs[14][20] ), .D(
        \regs[15][20] ), .S0(n1451), .S1(n1427), .Y(n1290) );
  MX4X1 U715 ( .A(\regs[28][21] ), .B(\regs[29][21] ), .C(\regs[30][21] ), .D(
        \regs[31][21] ), .S0(n1451), .S1(n1427), .Y(n1295) );
  MX4X1 U716 ( .A(\regs[12][21] ), .B(\regs[13][21] ), .C(\regs[14][21] ), .D(
        \regs[15][21] ), .S0(n1452), .S1(n1428), .Y(n1300) );
  MX4X1 U717 ( .A(\regs[28][22] ), .B(\regs[29][22] ), .C(\regs[30][22] ), .D(
        \regs[31][22] ), .S0(n1452), .S1(n1428), .Y(n1305) );
  MX4X1 U718 ( .A(\regs[12][22] ), .B(\regs[13][22] ), .C(\regs[14][22] ), .D(
        \regs[15][22] ), .S0(n1452), .S1(n1428), .Y(n1310) );
  MX4X1 U719 ( .A(\regs[28][23] ), .B(\regs[29][23] ), .C(\regs[30][23] ), .D(
        \regs[31][23] ), .S0(n1453), .S1(n1429), .Y(n1315) );
  MX4X1 U720 ( .A(\regs[12][23] ), .B(\regs[13][23] ), .C(\regs[14][23] ), .D(
        \regs[15][23] ), .S0(n1453), .S1(n1429), .Y(n1320) );
  MX4X1 U721 ( .A(\regs[28][24] ), .B(\regs[29][24] ), .C(\regs[30][24] ), .D(
        \regs[31][24] ), .S0(n1453), .S1(n1429), .Y(n1325) );
  MX4X1 U722 ( .A(\regs[12][24] ), .B(\regs[13][24] ), .C(\regs[14][24] ), .D(
        \regs[15][24] ), .S0(n1454), .S1(n1430), .Y(n1330) );
  MX4X1 U723 ( .A(\regs[28][25] ), .B(\regs[29][25] ), .C(\regs[30][25] ), .D(
        \regs[31][25] ), .S0(n1454), .S1(n1430), .Y(n1335) );
  MX4X1 U724 ( .A(\regs[12][25] ), .B(\regs[13][25] ), .C(\regs[14][25] ), .D(
        \regs[15][25] ), .S0(n1454), .S1(n1430), .Y(n1340) );
  MX4X1 U725 ( .A(\regs[28][26] ), .B(\regs[29][26] ), .C(\regs[30][26] ), .D(
        \regs[31][26] ), .S0(n1455), .S1(n1431), .Y(n1345) );
  MX4X1 U726 ( .A(\regs[12][26] ), .B(\regs[13][26] ), .C(\regs[14][26] ), .D(
        \regs[15][26] ), .S0(n1455), .S1(n1431), .Y(n1350) );
  MX4X1 U727 ( .A(\regs[28][27] ), .B(\regs[29][27] ), .C(\regs[30][27] ), .D(
        \regs[31][27] ), .S0(n1455), .S1(n1431), .Y(n1355) );
  MX4X1 U728 ( .A(\regs[12][27] ), .B(\regs[13][27] ), .C(\regs[14][27] ), .D(
        \regs[15][27] ), .S0(n1456), .S1(n1432), .Y(n1360) );
  MX4X1 U729 ( .A(\regs[28][28] ), .B(\regs[29][28] ), .C(\regs[30][28] ), .D(
        \regs[31][28] ), .S0(n1456), .S1(n1432), .Y(n1365) );
  MX4X1 U730 ( .A(\regs[12][28] ), .B(\regs[13][28] ), .C(\regs[14][28] ), .D(
        \regs[15][28] ), .S0(n1456), .S1(n1432), .Y(n1370) );
  MX4X1 U731 ( .A(\regs[28][29] ), .B(\regs[29][29] ), .C(\regs[30][29] ), .D(
        \regs[31][29] ), .S0(n1457), .S1(n1433), .Y(n1375) );
  MX4X1 U732 ( .A(\regs[12][29] ), .B(\regs[13][29] ), .C(\regs[14][29] ), .D(
        \regs[15][29] ), .S0(n1457), .S1(n1433), .Y(n1380) );
  MX4X1 U733 ( .A(\regs[28][30] ), .B(\regs[29][30] ), .C(\regs[30][30] ), .D(
        \regs[31][30] ), .S0(n1457), .S1(n1433), .Y(n1385) );
  MX4X1 U734 ( .A(\regs[12][30] ), .B(\regs[13][30] ), .C(\regs[14][30] ), .D(
        \regs[15][30] ), .S0(n1458), .S1(n1434), .Y(n1390) );
  MX4X1 U735 ( .A(\regs[28][31] ), .B(\regs[29][31] ), .C(\regs[30][31] ), .D(
        \regs[31][31] ), .S0(n1458), .S1(n1434), .Y(n1395) );
  MX4X1 U736 ( .A(\regs[12][31] ), .B(\regs[13][31] ), .C(\regs[14][31] ), .D(
        \regs[15][31] ), .S0(n1458), .S1(n1434), .Y(n1400) );
  MX4X1 U737 ( .A(\regs[24][26] ), .B(\regs[25][26] ), .C(\regs[26][26] ), .D(
        \regs[27][26] ), .S0(n1455), .S1(n1431), .Y(n1346) );
  MX4X1 U738 ( .A(\regs[8][26] ), .B(\regs[9][26] ), .C(\regs[10][26] ), .D(
        \regs[11][26] ), .S0(n1455), .S1(n1431), .Y(n1351) );
  MX4X1 U739 ( .A(\regs[24][27] ), .B(\regs[25][27] ), .C(\regs[26][27] ), .D(
        \regs[27][27] ), .S0(n1455), .S1(n1431), .Y(n1356) );
  MX4X1 U740 ( .A(\regs[8][27] ), .B(\regs[9][27] ), .C(\regs[10][27] ), .D(
        \regs[11][27] ), .S0(n1456), .S1(n1432), .Y(n1361) );
  MX4X1 U741 ( .A(\regs[24][28] ), .B(\regs[25][28] ), .C(\regs[26][28] ), .D(
        \regs[27][28] ), .S0(n1456), .S1(n1432), .Y(n1366) );
  MX4X1 U742 ( .A(\regs[8][28] ), .B(\regs[9][28] ), .C(\regs[10][28] ), .D(
        \regs[11][28] ), .S0(n1456), .S1(n1432), .Y(n1371) );
  MX4X1 U743 ( .A(\regs[24][29] ), .B(\regs[25][29] ), .C(\regs[26][29] ), .D(
        \regs[27][29] ), .S0(n1457), .S1(n1433), .Y(n1376) );
  MX4X1 U744 ( .A(\regs[8][29] ), .B(\regs[9][29] ), .C(\regs[10][29] ), .D(
        \regs[11][29] ), .S0(n1457), .S1(n1433), .Y(n1381) );
  MX4X1 U745 ( .A(n1833), .B(n1831), .C(n1832), .D(n1830), .S0(n2151), .S1(
        n2155), .Y(n1834) );
  MX4X1 U746 ( .A(\regs[16][0] ), .B(\regs[17][0] ), .C(\regs[18][0] ), .D(
        \regs[19][0] ), .S0(n2183), .S1(n2175), .Y(n1833) );
  MX4X1 U747 ( .A(\regs[24][0] ), .B(\regs[25][0] ), .C(\regs[26][0] ), .D(
        \regs[27][0] ), .S0(n2192), .S1(n2174), .Y(n1831) );
  MX4X1 U748 ( .A(\regs[20][0] ), .B(\regs[21][0] ), .C(\regs[22][0] ), .D(
        \regs[23][0] ), .S0(n2189), .S1(n2174), .Y(n1832) );
  MX4X1 U749 ( .A(n1843), .B(n1841), .C(n1842), .D(n1840), .S0(n2151), .S1(
        n2155), .Y(n1844) );
  MX4X1 U750 ( .A(\regs[16][1] ), .B(\regs[17][1] ), .C(\regs[18][1] ), .D(
        \regs[19][1] ), .S0(n2183), .S1(n2158), .Y(n1843) );
  MX4X1 U751 ( .A(\regs[24][1] ), .B(\regs[25][1] ), .C(\regs[26][1] ), .D(
        \regs[27][1] ), .S0(n2183), .S1(n2158), .Y(n1841) );
  MX4X1 U752 ( .A(\regs[20][1] ), .B(\regs[21][1] ), .C(\regs[22][1] ), .D(
        \regs[23][1] ), .S0(n2183), .S1(n2158), .Y(n1842) );
  MX4X1 U753 ( .A(n1853), .B(n1851), .C(n1852), .D(n1850), .S0(n2152), .S1(
        n2155), .Y(n1854) );
  MX4X1 U754 ( .A(\regs[16][2] ), .B(\regs[17][2] ), .C(\regs[18][2] ), .D(
        \regs[19][2] ), .S0(n2184), .S1(n2159), .Y(n1853) );
  MX4X1 U755 ( .A(\regs[24][2] ), .B(\regs[25][2] ), .C(\regs[26][2] ), .D(
        \regs[27][2] ), .S0(n2184), .S1(n2159), .Y(n1851) );
  MX4X1 U756 ( .A(\regs[20][2] ), .B(\regs[21][2] ), .C(\regs[22][2] ), .D(
        \regs[23][2] ), .S0(n2184), .S1(n2159), .Y(n1852) );
  MX4X1 U757 ( .A(n1863), .B(n1861), .C(n1862), .D(n1860), .S0(n2152), .S1(
        n2155), .Y(n1864) );
  MX4X1 U758 ( .A(\regs[16][3] ), .B(\regs[17][3] ), .C(\regs[18][3] ), .D(
        \regs[19][3] ), .S0(n2184), .S1(n2159), .Y(n1863) );
  MX4X1 U759 ( .A(\regs[24][3] ), .B(\regs[25][3] ), .C(\regs[26][3] ), .D(
        \regs[27][3] ), .S0(n2184), .S1(n2159), .Y(n1861) );
  MX4X1 U760 ( .A(\regs[20][3] ), .B(\regs[21][3] ), .C(\regs[22][3] ), .D(
        \regs[23][3] ), .S0(n2184), .S1(n2159), .Y(n1862) );
  MX4X1 U761 ( .A(n1873), .B(n1871), .C(n1872), .D(n1870), .S0(n2152), .S1(
        n2155), .Y(n1874) );
  MX4X1 U762 ( .A(\regs[16][4] ), .B(\regs[17][4] ), .C(\regs[18][4] ), .D(
        \regs[19][4] ), .S0(n2185), .S1(n2160), .Y(n1873) );
  MX4X1 U763 ( .A(\regs[24][4] ), .B(\regs[25][4] ), .C(\regs[26][4] ), .D(
        \regs[27][4] ), .S0(n2185), .S1(n2160), .Y(n1871) );
  MX4X1 U764 ( .A(\regs[20][4] ), .B(\regs[21][4] ), .C(\regs[22][4] ), .D(
        \regs[23][4] ), .S0(n2185), .S1(n2160), .Y(n1872) );
  MX4X1 U765 ( .A(n1883), .B(n1881), .C(n1882), .D(n1880), .S0(n2152), .S1(
        n2155), .Y(n1884) );
  MX4X1 U766 ( .A(\regs[16][5] ), .B(\regs[17][5] ), .C(\regs[18][5] ), .D(
        \regs[19][5] ), .S0(n2186), .S1(n2161), .Y(n1883) );
  MX4X1 U767 ( .A(\regs[24][5] ), .B(\regs[25][5] ), .C(\regs[26][5] ), .D(
        \regs[27][5] ), .S0(n2186), .S1(n2161), .Y(n1881) );
  MX4X1 U768 ( .A(\regs[20][5] ), .B(\regs[21][5] ), .C(\regs[22][5] ), .D(
        \regs[23][5] ), .S0(n2186), .S1(n2161), .Y(n1882) );
  MX4X1 U769 ( .A(n1893), .B(n1891), .C(n1892), .D(n1890), .S0(n2152), .S1(
        n2155), .Y(n1894) );
  MX4X1 U770 ( .A(\regs[16][6] ), .B(\regs[17][6] ), .C(\regs[18][6] ), .D(
        \regs[19][6] ), .S0(n2186), .S1(n2161), .Y(n1893) );
  MX4X1 U771 ( .A(\regs[24][6] ), .B(\regs[25][6] ), .C(\regs[26][6] ), .D(
        \regs[27][6] ), .S0(n2186), .S1(n2161), .Y(n1891) );
  MX4X1 U772 ( .A(\regs[20][6] ), .B(\regs[21][6] ), .C(\regs[22][6] ), .D(
        \regs[23][6] ), .S0(n2186), .S1(n2161), .Y(n1892) );
  MX4X1 U773 ( .A(n1903), .B(n1901), .C(n1902), .D(n1900), .S0(n2152), .S1(
        n2155), .Y(n1904) );
  MX4X1 U774 ( .A(\regs[16][7] ), .B(\regs[17][7] ), .C(\regs[18][7] ), .D(
        \regs[19][7] ), .S0(n2187), .S1(n2162), .Y(n1903) );
  MX4X1 U775 ( .A(\regs[24][7] ), .B(\regs[25][7] ), .C(\regs[26][7] ), .D(
        \regs[27][7] ), .S0(n2187), .S1(n2162), .Y(n1901) );
  MX4X1 U776 ( .A(\regs[20][7] ), .B(\regs[21][7] ), .C(\regs[22][7] ), .D(
        \regs[23][7] ), .S0(n2187), .S1(n2162), .Y(n1902) );
  MX4X1 U777 ( .A(n1913), .B(n1911), .C(n1912), .D(n1910), .S0(N25), .S1(n2155), .Y(n1914) );
  MX4X1 U778 ( .A(\regs[16][8] ), .B(\regs[17][8] ), .C(\regs[18][8] ), .D(
        \regs[19][8] ), .S0(n2188), .S1(n2163), .Y(n1913) );
  MX4X1 U779 ( .A(\regs[24][8] ), .B(\regs[25][8] ), .C(\regs[26][8] ), .D(
        \regs[27][8] ), .S0(n2188), .S1(n2163), .Y(n1911) );
  MX4X1 U780 ( .A(\regs[20][8] ), .B(\regs[21][8] ), .C(\regs[22][8] ), .D(
        \regs[23][8] ), .S0(n2188), .S1(n2163), .Y(n1912) );
  MX4X1 U781 ( .A(n1923), .B(n1921), .C(n1922), .D(n1920), .S0(n2153), .S1(N24), .Y(n1924) );
  MX4X1 U782 ( .A(\regs[16][9] ), .B(\regs[17][9] ), .C(\regs[18][9] ), .D(
        \regs[19][9] ), .S0(n2188), .S1(n2163), .Y(n1923) );
  MX4X1 U783 ( .A(\regs[24][9] ), .B(\regs[25][9] ), .C(\regs[26][9] ), .D(
        \regs[27][9] ), .S0(n2188), .S1(n2163), .Y(n1921) );
  MX4X1 U784 ( .A(\regs[20][9] ), .B(\regs[21][9] ), .C(\regs[22][9] ), .D(
        \regs[23][9] ), .S0(n2188), .S1(n2163), .Y(n1922) );
  MX4X1 U785 ( .A(n1933), .B(n1931), .C(n1932), .D(n1930), .S0(N25), .S1(n2155), .Y(n1934) );
  MX4X1 U786 ( .A(\regs[16][10] ), .B(\regs[17][10] ), .C(\regs[18][10] ), .D(
        \regs[19][10] ), .S0(n2189), .S1(n2164), .Y(n1933) );
  MX4X1 U787 ( .A(\regs[24][10] ), .B(\regs[25][10] ), .C(\regs[26][10] ), .D(
        \regs[27][10] ), .S0(n2189), .S1(n2164), .Y(n1931) );
  MX4X1 U788 ( .A(\regs[20][10] ), .B(\regs[21][10] ), .C(\regs[22][10] ), .D(
        \regs[23][10] ), .S0(n2189), .S1(n2164), .Y(n1932) );
  MX4X1 U789 ( .A(n1943), .B(n1941), .C(n1942), .D(n1940), .S0(n2152), .S1(
        n2155), .Y(n1944) );
  MX4X1 U790 ( .A(\regs[16][11] ), .B(\regs[17][11] ), .C(\regs[18][11] ), .D(
        \regs[19][11] ), .S0(n2190), .S1(n2165), .Y(n1943) );
  MX4X1 U791 ( .A(\regs[24][11] ), .B(\regs[25][11] ), .C(\regs[26][11] ), .D(
        \regs[27][11] ), .S0(n2190), .S1(n2165), .Y(n1941) );
  MX4X1 U792 ( .A(\regs[20][11] ), .B(\regs[21][11] ), .C(\regs[22][11] ), .D(
        \regs[23][11] ), .S0(n2190), .S1(n2165), .Y(n1942) );
  MX4X1 U793 ( .A(n1953), .B(n1951), .C(n1952), .D(n1950), .S0(n2152), .S1(
        n2155), .Y(n1954) );
  MX4X1 U794 ( .A(\regs[16][12] ), .B(\regs[17][12] ), .C(\regs[18][12] ), .D(
        \regs[19][12] ), .S0(n2190), .S1(n2165), .Y(n1953) );
  MX4X1 U795 ( .A(\regs[24][12] ), .B(\regs[25][12] ), .C(\regs[26][12] ), .D(
        \regs[27][12] ), .S0(n2190), .S1(n2165), .Y(n1951) );
  MX4X1 U796 ( .A(\regs[20][12] ), .B(\regs[21][12] ), .C(\regs[22][12] ), .D(
        \regs[23][12] ), .S0(n2190), .S1(n2165), .Y(n1952) );
  MX4X1 U797 ( .A(n1963), .B(n1961), .C(n1962), .D(n1960), .S0(N25), .S1(n2155), .Y(n1964) );
  MX4X1 U798 ( .A(\regs[16][13] ), .B(\regs[17][13] ), .C(\regs[18][13] ), .D(
        \regs[19][13] ), .S0(n2191), .S1(n2166), .Y(n1963) );
  MX4X1 U799 ( .A(\regs[24][13] ), .B(\regs[25][13] ), .C(\regs[26][13] ), .D(
        \regs[27][13] ), .S0(n2191), .S1(n2166), .Y(n1961) );
  MX4X1 U800 ( .A(\regs[20][13] ), .B(\regs[21][13] ), .C(\regs[22][13] ), .D(
        \regs[23][13] ), .S0(n2191), .S1(n2166), .Y(n1962) );
  MX4X1 U801 ( .A(n1973), .B(n1971), .C(n1972), .D(n1970), .S0(n2153), .S1(N24), .Y(n1974) );
  MX4X1 U802 ( .A(\regs[16][14] ), .B(\regs[17][14] ), .C(\regs[18][14] ), .D(
        \regs[19][14] ), .S0(n2192), .S1(n2167), .Y(n1973) );
  MX4X1 U803 ( .A(\regs[24][14] ), .B(\regs[25][14] ), .C(\regs[26][14] ), .D(
        \regs[27][14] ), .S0(n2192), .S1(n2167), .Y(n1971) );
  MX4X1 U804 ( .A(\regs[20][14] ), .B(\regs[21][14] ), .C(\regs[22][14] ), .D(
        \regs[23][14] ), .S0(n2192), .S1(n2167), .Y(n1972) );
  MX4X1 U805 ( .A(n1983), .B(n1981), .C(n1982), .D(n1980), .S0(n2153), .S1(
        n2155), .Y(n1984) );
  MX4X1 U806 ( .A(\regs[16][15] ), .B(\regs[17][15] ), .C(\regs[18][15] ), .D(
        \regs[19][15] ), .S0(n2192), .S1(n2167), .Y(n1983) );
  MX4X1 U807 ( .A(\regs[24][15] ), .B(\regs[25][15] ), .C(\regs[26][15] ), .D(
        \regs[27][15] ), .S0(n2192), .S1(n2167), .Y(n1981) );
  MX4X1 U808 ( .A(\regs[20][15] ), .B(\regs[21][15] ), .C(\regs[22][15] ), .D(
        \regs[23][15] ), .S0(n2192), .S1(n2167), .Y(n1982) );
  MX4X1 U809 ( .A(n1993), .B(n1991), .C(n1992), .D(n1990), .S0(n2153), .S1(N24), .Y(n1994) );
  MX4X1 U810 ( .A(\regs[16][16] ), .B(\regs[17][16] ), .C(\regs[18][16] ), .D(
        \regs[19][16] ), .S0(n2193), .S1(n2168), .Y(n1993) );
  MX4X1 U811 ( .A(\regs[24][16] ), .B(\regs[25][16] ), .C(\regs[26][16] ), .D(
        \regs[27][16] ), .S0(n2193), .S1(n2168), .Y(n1991) );
  MX4X1 U812 ( .A(\regs[20][16] ), .B(\regs[21][16] ), .C(\regs[22][16] ), .D(
        \regs[23][16] ), .S0(n2193), .S1(n2168), .Y(n1992) );
  MX4X1 U813 ( .A(n2003), .B(n2001), .C(n2002), .D(n2000), .S0(n2153), .S1(N24), .Y(n2004) );
  MX4X1 U814 ( .A(\regs[16][17] ), .B(\regs[17][17] ), .C(\regs[18][17] ), .D(
        \regs[19][17] ), .S0(n2194), .S1(n2169), .Y(n2003) );
  MX4X1 U815 ( .A(\regs[24][17] ), .B(\regs[25][17] ), .C(\regs[26][17] ), .D(
        \regs[27][17] ), .S0(n2194), .S1(n2169), .Y(n2001) );
  MX4X1 U816 ( .A(\regs[20][17] ), .B(\regs[21][17] ), .C(\regs[22][17] ), .D(
        \regs[23][17] ), .S0(n2194), .S1(n2169), .Y(n2002) );
  MX4X1 U817 ( .A(n2013), .B(n2011), .C(n2012), .D(n2010), .S0(n2153), .S1(N24), .Y(n2014) );
  MX4X1 U818 ( .A(\regs[16][18] ), .B(\regs[17][18] ), .C(\regs[18][18] ), .D(
        \regs[19][18] ), .S0(n2194), .S1(n2169), .Y(n2013) );
  MX4X1 U819 ( .A(\regs[24][18] ), .B(\regs[25][18] ), .C(\regs[26][18] ), .D(
        \regs[27][18] ), .S0(n2194), .S1(n2169), .Y(n2011) );
  MX4X1 U820 ( .A(\regs[20][18] ), .B(\regs[21][18] ), .C(\regs[22][18] ), .D(
        \regs[23][18] ), .S0(n2194), .S1(n2169), .Y(n2012) );
  MX4X1 U821 ( .A(n2023), .B(n2021), .C(n2022), .D(n2020), .S0(n2153), .S1(N24), .Y(n2024) );
  MX4X1 U822 ( .A(\regs[16][19] ), .B(\regs[17][19] ), .C(\regs[18][19] ), .D(
        \regs[19][19] ), .S0(n2195), .S1(n2170), .Y(n2023) );
  MX4X1 U823 ( .A(\regs[24][19] ), .B(\regs[25][19] ), .C(\regs[26][19] ), .D(
        \regs[27][19] ), .S0(n2195), .S1(n2170), .Y(n2021) );
  MX4X1 U824 ( .A(\regs[20][19] ), .B(\regs[21][19] ), .C(\regs[22][19] ), .D(
        \regs[23][19] ), .S0(n2195), .S1(n2170), .Y(n2022) );
  MX4X1 U825 ( .A(n2033), .B(n2031), .C(n2032), .D(n2030), .S0(n2153), .S1(N24), .Y(n2034) );
  MX4X1 U826 ( .A(\regs[16][20] ), .B(\regs[17][20] ), .C(\regs[18][20] ), .D(
        \regs[19][20] ), .S0(n2196), .S1(n2171), .Y(n2033) );
  MX4X1 U827 ( .A(\regs[24][20] ), .B(\regs[25][20] ), .C(\regs[26][20] ), .D(
        \regs[27][20] ), .S0(n2196), .S1(n2171), .Y(n2031) );
  MX4X1 U828 ( .A(\regs[20][20] ), .B(\regs[21][20] ), .C(\regs[22][20] ), .D(
        \regs[23][20] ), .S0(n2196), .S1(n2171), .Y(n2032) );
  MX4X1 U829 ( .A(n2043), .B(n2041), .C(n2042), .D(n2040), .S0(N25), .S1(N24), 
        .Y(n2044) );
  MX4X1 U830 ( .A(\regs[16][21] ), .B(\regs[17][21] ), .C(\regs[18][21] ), .D(
        \regs[19][21] ), .S0(n2196), .S1(n2171), .Y(n2043) );
  MX4X1 U831 ( .A(\regs[24][21] ), .B(\regs[25][21] ), .C(\regs[26][21] ), .D(
        \regs[27][21] ), .S0(n2196), .S1(n2171), .Y(n2041) );
  MX4X1 U832 ( .A(\regs[20][21] ), .B(\regs[21][21] ), .C(\regs[22][21] ), .D(
        \regs[23][21] ), .S0(n2196), .S1(n2171), .Y(n2042) );
  MX4X1 U833 ( .A(n2053), .B(n2051), .C(n2052), .D(n2050), .S0(N25), .S1(N24), 
        .Y(n2054) );
  MX4X1 U834 ( .A(\regs[16][22] ), .B(\regs[17][22] ), .C(\regs[18][22] ), .D(
        \regs[19][22] ), .S0(n2197), .S1(n2172), .Y(n2053) );
  MX4X1 U835 ( .A(\regs[24][22] ), .B(\regs[25][22] ), .C(\regs[26][22] ), .D(
        \regs[27][22] ), .S0(n2197), .S1(n2172), .Y(n2051) );
  MX4X1 U836 ( .A(\regs[20][22] ), .B(\regs[21][22] ), .C(\regs[22][22] ), .D(
        \regs[23][22] ), .S0(n2197), .S1(n2172), .Y(n2052) );
  MX4X1 U837 ( .A(n2063), .B(n2061), .C(n2062), .D(n2060), .S0(n2151), .S1(N24), .Y(n2064) );
  MX4X1 U838 ( .A(\regs[16][23] ), .B(\regs[17][23] ), .C(\regs[18][23] ), .D(
        \regs[19][23] ), .S0(n2198), .S1(n2173), .Y(n2063) );
  MX4X1 U839 ( .A(\regs[24][23] ), .B(\regs[25][23] ), .C(\regs[26][23] ), .D(
        \regs[27][23] ), .S0(n2198), .S1(n2173), .Y(n2061) );
  MX4X1 U840 ( .A(\regs[20][23] ), .B(\regs[21][23] ), .C(\regs[22][23] ), .D(
        \regs[23][23] ), .S0(n2198), .S1(n2173), .Y(n2062) );
  MX4X1 U841 ( .A(n2073), .B(n2071), .C(n2072), .D(n2070), .S0(n2152), .S1(
        n2155), .Y(n2074) );
  MX4X1 U842 ( .A(\regs[16][24] ), .B(\regs[17][24] ), .C(\regs[18][24] ), .D(
        \regs[19][24] ), .S0(n2198), .S1(n2173), .Y(n2073) );
  MX4X1 U843 ( .A(\regs[24][24] ), .B(\regs[25][24] ), .C(\regs[26][24] ), .D(
        \regs[27][24] ), .S0(n2198), .S1(n2173), .Y(n2071) );
  MX4X1 U844 ( .A(\regs[20][24] ), .B(\regs[21][24] ), .C(\regs[22][24] ), .D(
        \regs[23][24] ), .S0(n2198), .S1(n2173), .Y(n2072) );
  MX4X1 U845 ( .A(n2083), .B(n2081), .C(n2082), .D(n2080), .S0(N25), .S1(N24), 
        .Y(n2084) );
  MX4X1 U846 ( .A(\regs[16][25] ), .B(\regs[17][25] ), .C(\regs[18][25] ), .D(
        \regs[19][25] ), .S0(n2199), .S1(n2174), .Y(n2083) );
  MX4X1 U847 ( .A(\regs[24][25] ), .B(\regs[25][25] ), .C(\regs[26][25] ), .D(
        \regs[27][25] ), .S0(n2199), .S1(n2174), .Y(n2081) );
  MX4X1 U848 ( .A(\regs[20][25] ), .B(\regs[21][25] ), .C(\regs[22][25] ), .D(
        \regs[23][25] ), .S0(n2199), .S1(n2174), .Y(n2082) );
  MX4X1 U849 ( .A(n2093), .B(n2091), .C(n2092), .D(n2090), .S0(n2152), .S1(N24), .Y(n2094) );
  MX4X1 U850 ( .A(\regs[16][26] ), .B(\regs[17][26] ), .C(\regs[18][26] ), .D(
        \regs[19][26] ), .S0(n2200), .S1(n2175), .Y(n2093) );
  MX4X1 U851 ( .A(\regs[24][26] ), .B(\regs[25][26] ), .C(\regs[26][26] ), .D(
        \regs[27][26] ), .S0(n2200), .S1(n2175), .Y(n2091) );
  MX4X1 U852 ( .A(\regs[20][26] ), .B(\regs[21][26] ), .C(\regs[22][26] ), .D(
        \regs[23][26] ), .S0(n2200), .S1(n2175), .Y(n2092) );
  MX4X1 U853 ( .A(n2103), .B(n2101), .C(n2102), .D(n2100), .S0(n2151), .S1(N24), .Y(n2104) );
  MX4X1 U854 ( .A(\regs[16][27] ), .B(\regs[17][27] ), .C(\regs[18][27] ), .D(
        \regs[19][27] ), .S0(n2200), .S1(n2175), .Y(n2103) );
  MX4X1 U855 ( .A(\regs[24][27] ), .B(\regs[25][27] ), .C(\regs[26][27] ), .D(
        \regs[27][27] ), .S0(n2200), .S1(n2175), .Y(n2101) );
  MX4X1 U856 ( .A(\regs[20][27] ), .B(\regs[21][27] ), .C(\regs[22][27] ), .D(
        \regs[23][27] ), .S0(n2200), .S1(n2175), .Y(n2102) );
  MX4X1 U857 ( .A(n2113), .B(n2111), .C(n2112), .D(n2110), .S0(n2151), .S1(N24), .Y(n2114) );
  MX4X1 U858 ( .A(\regs[16][28] ), .B(\regs[17][28] ), .C(\regs[18][28] ), .D(
        \regs[19][28] ), .S0(n2201), .S1(n2176), .Y(n2113) );
  MX4X1 U859 ( .A(\regs[24][28] ), .B(\regs[25][28] ), .C(\regs[26][28] ), .D(
        \regs[27][28] ), .S0(n2201), .S1(n2176), .Y(n2111) );
  MX4X1 U860 ( .A(\regs[20][28] ), .B(\regs[21][28] ), .C(\regs[22][28] ), .D(
        \regs[23][28] ), .S0(n2201), .S1(n2176), .Y(n2112) );
  MX4X1 U861 ( .A(n2123), .B(n2121), .C(n2122), .D(n2120), .S0(n2151), .S1(N24), .Y(n2124) );
  MX4X1 U862 ( .A(\regs[16][29] ), .B(\regs[17][29] ), .C(\regs[18][29] ), .D(
        \regs[19][29] ), .S0(n2202), .S1(n2177), .Y(n2123) );
  MX4X1 U863 ( .A(\regs[24][29] ), .B(\regs[25][29] ), .C(\regs[26][29] ), .D(
        \regs[27][29] ), .S0(n2202), .S1(n2177), .Y(n2121) );
  MX4X1 U864 ( .A(\regs[20][29] ), .B(\regs[21][29] ), .C(\regs[22][29] ), .D(
        \regs[23][29] ), .S0(n2202), .S1(n2177), .Y(n2122) );
  MX4X1 U865 ( .A(n2133), .B(n2131), .C(n2132), .D(n2130), .S0(n2151), .S1(
        n2155), .Y(n2134) );
  MX4X1 U866 ( .A(\regs[16][30] ), .B(\regs[17][30] ), .C(\regs[18][30] ), .D(
        \regs[19][30] ), .S0(n2202), .S1(n2177), .Y(n2133) );
  MX4X1 U867 ( .A(\regs[24][30] ), .B(\regs[25][30] ), .C(\regs[26][30] ), .D(
        \regs[27][30] ), .S0(n2202), .S1(n2177), .Y(n2131) );
  MX4X1 U868 ( .A(\regs[20][30] ), .B(\regs[21][30] ), .C(\regs[22][30] ), .D(
        \regs[23][30] ), .S0(n2202), .S1(n2177), .Y(n2132) );
  MX4X1 U869 ( .A(n2143), .B(n2141), .C(n2142), .D(n2140), .S0(n2151), .S1(N24), .Y(n2144) );
  MX4X1 U870 ( .A(\regs[16][31] ), .B(\regs[17][31] ), .C(\regs[18][31] ), .D(
        \regs[19][31] ), .S0(n2203), .S1(n2178), .Y(n2143) );
  MX4X1 U871 ( .A(\regs[24][31] ), .B(\regs[25][31] ), .C(\regs[26][31] ), .D(
        \regs[27][31] ), .S0(n2203), .S1(n2178), .Y(n2141) );
  MX4X1 U872 ( .A(\regs[20][31] ), .B(\regs[21][31] ), .C(\regs[22][31] ), .D(
        \regs[23][31] ), .S0(n2203), .S1(n2178), .Y(n2142) );
  MX4X1 U873 ( .A(n49), .B(n47), .C(n48), .D(n45), .S0(n1407), .S1(n1410), .Y(
        n51) );
  MX4X1 U874 ( .A(\regs[16][0] ), .B(\regs[17][0] ), .C(\regs[18][0] ), .D(
        \regs[19][0] ), .S0(n1438), .S1(n1423), .Y(n49) );
  MX4X1 U875 ( .A(\regs[24][0] ), .B(\regs[25][0] ), .C(\regs[26][0] ), .D(
        \regs[27][0] ), .S0(n1444), .S1(n1419), .Y(n47) );
  MX4X1 U876 ( .A(\regs[20][0] ), .B(\regs[21][0] ), .C(\regs[22][0] ), .D(
        \regs[23][0] ), .S0(n1447), .S1(n1422), .Y(n48) );
  MX4X1 U877 ( .A(n69), .B(n63), .C(n65), .D(n60), .S0(n1406), .S1(n1410), .Y(
        n71) );
  MX4X1 U878 ( .A(\regs[16][1] ), .B(\regs[17][1] ), .C(\regs[18][1] ), .D(
        \regs[19][1] ), .S0(n1438), .S1(n1414), .Y(n69) );
  MX4X1 U879 ( .A(\regs[24][1] ), .B(\regs[25][1] ), .C(\regs[26][1] ), .D(
        \regs[27][1] ), .S0(n1438), .S1(n1414), .Y(n63) );
  MX4X1 U880 ( .A(\regs[20][1] ), .B(\regs[21][1] ), .C(\regs[22][1] ), .D(
        \regs[23][1] ), .S0(n1438), .S1(n1414), .Y(n65) );
  MX4X1 U881 ( .A(n84), .B(n80), .C(n82), .D(n79), .S0(n1406), .S1(n1410), .Y(
        n85) );
  MX4X1 U882 ( .A(\regs[16][2] ), .B(\regs[17][2] ), .C(\regs[18][2] ), .D(
        \regs[19][2] ), .S0(n1439), .S1(n1415), .Y(n84) );
  MX4X1 U883 ( .A(\regs[24][2] ), .B(\regs[25][2] ), .C(\regs[26][2] ), .D(
        \regs[27][2] ), .S0(n1439), .S1(n1415), .Y(n80) );
  MX4X1 U884 ( .A(\regs[20][2] ), .B(\regs[21][2] ), .C(\regs[22][2] ), .D(
        \regs[23][2] ), .S0(n1439), .S1(n1415), .Y(n82) );
  MX4X1 U885 ( .A(n1118), .B(n1116), .C(n1117), .D(n1115), .S0(n1406), .S1(
        n1410), .Y(n1119) );
  MX4X1 U886 ( .A(\regs[16][3] ), .B(\regs[17][3] ), .C(\regs[18][3] ), .D(
        \regs[19][3] ), .S0(n1439), .S1(n1415), .Y(n1118) );
  MX4X1 U887 ( .A(\regs[24][3] ), .B(\regs[25][3] ), .C(\regs[26][3] ), .D(
        \regs[27][3] ), .S0(n1439), .S1(n1415), .Y(n1116) );
  MX4X1 U888 ( .A(\regs[20][3] ), .B(\regs[21][3] ), .C(\regs[22][3] ), .D(
        \regs[23][3] ), .S0(n1439), .S1(n1415), .Y(n1117) );
  MX4X1 U889 ( .A(n1128), .B(n1126), .C(n1127), .D(n1125), .S0(n1406), .S1(
        n1410), .Y(n1129) );
  MX4X1 U890 ( .A(\regs[16][4] ), .B(\regs[17][4] ), .C(\regs[18][4] ), .D(
        \regs[19][4] ), .S0(n1440), .S1(n1416), .Y(n1128) );
  MX4X1 U891 ( .A(\regs[24][4] ), .B(\regs[25][4] ), .C(\regs[26][4] ), .D(
        \regs[27][4] ), .S0(n1440), .S1(n1416), .Y(n1126) );
  MX4X1 U892 ( .A(\regs[20][4] ), .B(\regs[21][4] ), .C(\regs[22][4] ), .D(
        \regs[23][4] ), .S0(n1440), .S1(n1416), .Y(n1127) );
  MX4X1 U893 ( .A(n1138), .B(n1136), .C(n1137), .D(n1135), .S0(n1406), .S1(
        n1410), .Y(n1139) );
  MX4X1 U894 ( .A(\regs[16][5] ), .B(\regs[17][5] ), .C(\regs[18][5] ), .D(
        \regs[19][5] ), .S0(n1441), .S1(n1417), .Y(n1138) );
  MX4X1 U895 ( .A(\regs[24][5] ), .B(\regs[25][5] ), .C(\regs[26][5] ), .D(
        \regs[27][5] ), .S0(n1441), .S1(n1417), .Y(n1136) );
  MX4X1 U896 ( .A(\regs[20][5] ), .B(\regs[21][5] ), .C(\regs[22][5] ), .D(
        \regs[23][5] ), .S0(n1441), .S1(n1417), .Y(n1137) );
  MX4X1 U897 ( .A(n1148), .B(n1146), .C(n1147), .D(n1145), .S0(n1406), .S1(
        n1410), .Y(n1149) );
  MX4X1 U898 ( .A(\regs[16][6] ), .B(\regs[17][6] ), .C(\regs[18][6] ), .D(
        \regs[19][6] ), .S0(n1441), .S1(n1417), .Y(n1148) );
  MX4X1 U899 ( .A(\regs[24][6] ), .B(\regs[25][6] ), .C(\regs[26][6] ), .D(
        \regs[27][6] ), .S0(n1441), .S1(n1417), .Y(n1146) );
  MX4X1 U900 ( .A(\regs[20][6] ), .B(\regs[21][6] ), .C(\regs[22][6] ), .D(
        \regs[23][6] ), .S0(n1441), .S1(n1417), .Y(n1147) );
  MX4X1 U901 ( .A(n1158), .B(n1156), .C(n1157), .D(n1155), .S0(n1406), .S1(
        n1410), .Y(n1159) );
  MX4X1 U902 ( .A(\regs[16][7] ), .B(\regs[17][7] ), .C(\regs[18][7] ), .D(
        \regs[19][7] ), .S0(n1442), .S1(n1418), .Y(n1158) );
  MX4X1 U903 ( .A(\regs[24][7] ), .B(\regs[25][7] ), .C(\regs[26][7] ), .D(
        \regs[27][7] ), .S0(n1442), .S1(n1418), .Y(n1156) );
  MX4X1 U904 ( .A(\regs[20][7] ), .B(\regs[21][7] ), .C(\regs[22][7] ), .D(
        \regs[23][7] ), .S0(n1442), .S1(n1418), .Y(n1157) );
  MX4X1 U905 ( .A(n1168), .B(n1166), .C(n1167), .D(n1165), .S0(N15), .S1(n1410), .Y(n1169) );
  MX4X1 U906 ( .A(\regs[16][8] ), .B(\regs[17][8] ), .C(\regs[18][8] ), .D(
        \regs[19][8] ), .S0(n1443), .S1(n1419), .Y(n1168) );
  MX4X1 U907 ( .A(\regs[24][8] ), .B(\regs[25][8] ), .C(\regs[26][8] ), .D(
        \regs[27][8] ), .S0(n1443), .S1(n1419), .Y(n1166) );
  MX4X1 U908 ( .A(\regs[20][8] ), .B(\regs[21][8] ), .C(\regs[22][8] ), .D(
        \regs[23][8] ), .S0(n1443), .S1(n1419), .Y(n1167) );
  MX4X1 U909 ( .A(n1178), .B(n1176), .C(n1177), .D(n1175), .S0(N15), .S1(n1410), .Y(n1179) );
  MX4X1 U910 ( .A(\regs[16][9] ), .B(\regs[17][9] ), .C(\regs[18][9] ), .D(
        \regs[19][9] ), .S0(n1443), .S1(n1419), .Y(n1178) );
  MX4X1 U911 ( .A(\regs[24][9] ), .B(\regs[25][9] ), .C(\regs[26][9] ), .D(
        \regs[27][9] ), .S0(n1443), .S1(n1419), .Y(n1176) );
  MX4X1 U912 ( .A(\regs[20][9] ), .B(\regs[21][9] ), .C(\regs[22][9] ), .D(
        \regs[23][9] ), .S0(n1443), .S1(n1419), .Y(n1177) );
  MX4X1 U913 ( .A(n1188), .B(n1186), .C(n1187), .D(n1185), .S0(N15), .S1(n1410), .Y(n1189) );
  MX4X1 U914 ( .A(\regs[16][10] ), .B(\regs[17][10] ), .C(\regs[18][10] ), .D(
        \regs[19][10] ), .S0(n1444), .S1(n1420), .Y(n1188) );
  MX4X1 U915 ( .A(\regs[24][10] ), .B(\regs[25][10] ), .C(\regs[26][10] ), .D(
        \regs[27][10] ), .S0(n1444), .S1(n1420), .Y(n1186) );
  MX4X1 U916 ( .A(\regs[20][10] ), .B(\regs[21][10] ), .C(\regs[22][10] ), .D(
        \regs[23][10] ), .S0(n1444), .S1(n1420), .Y(n1187) );
  MX4X1 U917 ( .A(n1198), .B(n1196), .C(n1197), .D(n1195), .S0(n1408), .S1(
        n1410), .Y(n1199) );
  MX4X1 U918 ( .A(\regs[16][11] ), .B(\regs[17][11] ), .C(\regs[18][11] ), .D(
        \regs[19][11] ), .S0(n1445), .S1(n1421), .Y(n1198) );
  MX4X1 U919 ( .A(\regs[24][11] ), .B(\regs[25][11] ), .C(\regs[26][11] ), .D(
        \regs[27][11] ), .S0(n1445), .S1(n1421), .Y(n1196) );
  MX4X1 U920 ( .A(\regs[20][11] ), .B(\regs[21][11] ), .C(\regs[22][11] ), .D(
        \regs[23][11] ), .S0(n1445), .S1(n1421), .Y(n1197) );
  MX4X1 U921 ( .A(n1208), .B(n1206), .C(n1207), .D(n1205), .S0(n1406), .S1(
        n1410), .Y(n1209) );
  MX4X1 U922 ( .A(\regs[16][12] ), .B(\regs[17][12] ), .C(\regs[18][12] ), .D(
        \regs[19][12] ), .S0(n1445), .S1(n1421), .Y(n1208) );
  MX4X1 U923 ( .A(\regs[24][12] ), .B(\regs[25][12] ), .C(\regs[26][12] ), .D(
        \regs[27][12] ), .S0(n1445), .S1(n1421), .Y(n1206) );
  MX4X1 U924 ( .A(\regs[20][12] ), .B(\regs[21][12] ), .C(\regs[22][12] ), .D(
        \regs[23][12] ), .S0(n1445), .S1(n1421), .Y(n1207) );
  MX4X1 U925 ( .A(n1218), .B(n1216), .C(n1217), .D(n1215), .S0(n1408), .S1(
        n1410), .Y(n1219) );
  MX4X1 U926 ( .A(\regs[16][13] ), .B(\regs[17][13] ), .C(\regs[18][13] ), .D(
        \regs[19][13] ), .S0(n1446), .S1(n1422), .Y(n1218) );
  MX4X1 U927 ( .A(\regs[24][13] ), .B(\regs[25][13] ), .C(\regs[26][13] ), .D(
        \regs[27][13] ), .S0(n1446), .S1(n1422), .Y(n1216) );
  MX4X1 U928 ( .A(\regs[20][13] ), .B(\regs[21][13] ), .C(\regs[22][13] ), .D(
        \regs[23][13] ), .S0(n1446), .S1(n1422), .Y(n1217) );
  MX4X1 U929 ( .A(n1228), .B(n1226), .C(n1227), .D(n1225), .S0(n1407), .S1(N14), .Y(n1229) );
  MX4X1 U930 ( .A(\regs[16][14] ), .B(\regs[17][14] ), .C(\regs[18][14] ), .D(
        \regs[19][14] ), .S0(n1447), .S1(n1423), .Y(n1228) );
  MX4X1 U931 ( .A(\regs[24][14] ), .B(\regs[25][14] ), .C(\regs[26][14] ), .D(
        \regs[27][14] ), .S0(n1447), .S1(n1423), .Y(n1226) );
  MX4X1 U932 ( .A(\regs[20][14] ), .B(\regs[21][14] ), .C(\regs[22][14] ), .D(
        \regs[23][14] ), .S0(n1447), .S1(n1423), .Y(n1227) );
  MX4X1 U933 ( .A(n1238), .B(n1236), .C(n1237), .D(n1235), .S0(n1407), .S1(
        n1410), .Y(n1239) );
  MX4X1 U934 ( .A(\regs[16][15] ), .B(\regs[17][15] ), .C(\regs[18][15] ), .D(
        \regs[19][15] ), .S0(n1447), .S1(n1423), .Y(n1238) );
  MX4X1 U935 ( .A(\regs[24][15] ), .B(\regs[25][15] ), .C(\regs[26][15] ), .D(
        \regs[27][15] ), .S0(n1447), .S1(n1423), .Y(n1236) );
  MX4X1 U936 ( .A(\regs[20][15] ), .B(\regs[21][15] ), .C(\regs[22][15] ), .D(
        \regs[23][15] ), .S0(n1447), .S1(n1423), .Y(n1237) );
  MX4X1 U937 ( .A(n1248), .B(n1246), .C(n1247), .D(n1245), .S0(n1407), .S1(N14), .Y(n1249) );
  MX4X1 U938 ( .A(\regs[16][16] ), .B(\regs[17][16] ), .C(\regs[18][16] ), .D(
        \regs[19][16] ), .S0(n1448), .S1(n1424), .Y(n1248) );
  MX4X1 U939 ( .A(\regs[24][16] ), .B(\regs[25][16] ), .C(\regs[26][16] ), .D(
        \regs[27][16] ), .S0(n1448), .S1(n1424), .Y(n1246) );
  MX4X1 U940 ( .A(\regs[20][16] ), .B(\regs[21][16] ), .C(\regs[22][16] ), .D(
        \regs[23][16] ), .S0(n1448), .S1(n1424), .Y(n1247) );
  MX4X1 U941 ( .A(n1258), .B(n1256), .C(n1257), .D(n1255), .S0(n1407), .S1(N14), .Y(n1259) );
  MX4X1 U942 ( .A(\regs[16][17] ), .B(\regs[17][17] ), .C(\regs[18][17] ), .D(
        \regs[19][17] ), .S0(n1449), .S1(n1425), .Y(n1258) );
  MX4X1 U943 ( .A(\regs[24][17] ), .B(\regs[25][17] ), .C(\regs[26][17] ), .D(
        \regs[27][17] ), .S0(n1449), .S1(n1425), .Y(n1256) );
  MX4X1 U944 ( .A(\regs[20][17] ), .B(\regs[21][17] ), .C(\regs[22][17] ), .D(
        \regs[23][17] ), .S0(n1449), .S1(n1425), .Y(n1257) );
  MX4X1 U945 ( .A(n1268), .B(n1266), .C(n1267), .D(n1265), .S0(n1407), .S1(N14), .Y(n1269) );
  MX4X1 U946 ( .A(\regs[16][18] ), .B(\regs[17][18] ), .C(\regs[18][18] ), .D(
        \regs[19][18] ), .S0(n1449), .S1(n1425), .Y(n1268) );
  MX4X1 U947 ( .A(\regs[24][18] ), .B(\regs[25][18] ), .C(\regs[26][18] ), .D(
        \regs[27][18] ), .S0(n1449), .S1(n1425), .Y(n1266) );
  MX4X1 U948 ( .A(\regs[20][18] ), .B(\regs[21][18] ), .C(\regs[22][18] ), .D(
        \regs[23][18] ), .S0(n1449), .S1(n1425), .Y(n1267) );
  MX4X1 U949 ( .A(n1278), .B(n1276), .C(n1277), .D(n1275), .S0(n1407), .S1(N14), .Y(n1279) );
  MX4X1 U950 ( .A(\regs[16][19] ), .B(\regs[17][19] ), .C(\regs[18][19] ), .D(
        \regs[19][19] ), .S0(n1450), .S1(n1426), .Y(n1278) );
  MX4X1 U951 ( .A(\regs[24][19] ), .B(\regs[25][19] ), .C(\regs[26][19] ), .D(
        \regs[27][19] ), .S0(n1450), .S1(n1426), .Y(n1276) );
  MX4X1 U952 ( .A(\regs[20][19] ), .B(\regs[21][19] ), .C(\regs[22][19] ), .D(
        \regs[23][19] ), .S0(n1450), .S1(n1426), .Y(n1277) );
  MX4X1 U953 ( .A(n1288), .B(n1286), .C(n1287), .D(n1285), .S0(n1407), .S1(N14), .Y(n1289) );
  MX4X1 U954 ( .A(\regs[16][20] ), .B(\regs[17][20] ), .C(\regs[18][20] ), .D(
        \regs[19][20] ), .S0(n1451), .S1(n1427), .Y(n1288) );
  MX4X1 U955 ( .A(\regs[24][20] ), .B(\regs[25][20] ), .C(\regs[26][20] ), .D(
        \regs[27][20] ), .S0(n1451), .S1(n1427), .Y(n1286) );
  MX4X1 U956 ( .A(\regs[20][20] ), .B(\regs[21][20] ), .C(\regs[22][20] ), .D(
        \regs[23][20] ), .S0(n1451), .S1(n1427), .Y(n1287) );
  MX4X1 U957 ( .A(n1298), .B(n1296), .C(n1297), .D(n1295), .S0(N15), .S1(N14), 
        .Y(n1299) );
  MX4X1 U958 ( .A(\regs[16][21] ), .B(\regs[17][21] ), .C(\regs[18][21] ), .D(
        \regs[19][21] ), .S0(n1451), .S1(n1427), .Y(n1298) );
  MX4X1 U959 ( .A(\regs[24][21] ), .B(\regs[25][21] ), .C(\regs[26][21] ), .D(
        \regs[27][21] ), .S0(n1451), .S1(n1427), .Y(n1296) );
  MX4X1 U960 ( .A(\regs[20][21] ), .B(\regs[21][21] ), .C(\regs[22][21] ), .D(
        \regs[23][21] ), .S0(n1451), .S1(n1427), .Y(n1297) );
  MX4X1 U961 ( .A(n1308), .B(n1306), .C(n1307), .D(n1305), .S0(N15), .S1(N14), 
        .Y(n1309) );
  MX4X1 U962 ( .A(\regs[16][22] ), .B(\regs[17][22] ), .C(\regs[18][22] ), .D(
        \regs[19][22] ), .S0(n1452), .S1(n1428), .Y(n1308) );
  MX4X1 U963 ( .A(\regs[24][22] ), .B(\regs[25][22] ), .C(\regs[26][22] ), .D(
        \regs[27][22] ), .S0(n1452), .S1(n1428), .Y(n1306) );
  MX4X1 U964 ( .A(\regs[20][22] ), .B(\regs[21][22] ), .C(\regs[22][22] ), .D(
        \regs[23][22] ), .S0(n1452), .S1(n1428), .Y(n1307) );
  MX4X1 U965 ( .A(n1318), .B(n1316), .C(n1317), .D(n1315), .S0(N15), .S1(N14), 
        .Y(n1319) );
  MX4X1 U966 ( .A(\regs[16][23] ), .B(\regs[17][23] ), .C(\regs[18][23] ), .D(
        \regs[19][23] ), .S0(n1453), .S1(n1429), .Y(n1318) );
  MX4X1 U967 ( .A(\regs[24][23] ), .B(\regs[25][23] ), .C(\regs[26][23] ), .D(
        \regs[27][23] ), .S0(n1453), .S1(n1429), .Y(n1316) );
  MX4X1 U968 ( .A(\regs[20][23] ), .B(\regs[21][23] ), .C(\regs[22][23] ), .D(
        \regs[23][23] ), .S0(n1453), .S1(n1429), .Y(n1317) );
  MX4X1 U969 ( .A(n1328), .B(n1326), .C(n1327), .D(n1325), .S0(n1408), .S1(
        n1410), .Y(n1329) );
  MX4X1 U970 ( .A(\regs[16][24] ), .B(\regs[17][24] ), .C(\regs[18][24] ), .D(
        \regs[19][24] ), .S0(n1453), .S1(n1429), .Y(n1328) );
  MX4X1 U971 ( .A(\regs[24][24] ), .B(\regs[25][24] ), .C(\regs[26][24] ), .D(
        \regs[27][24] ), .S0(n1453), .S1(n1429), .Y(n1326) );
  MX4X1 U972 ( .A(\regs[20][24] ), .B(\regs[21][24] ), .C(\regs[22][24] ), .D(
        \regs[23][24] ), .S0(n1453), .S1(n1429), .Y(n1327) );
  MX4X1 U973 ( .A(n1338), .B(n1336), .C(n1337), .D(n1335), .S0(N15), .S1(N14), 
        .Y(n1339) );
  MX4X1 U974 ( .A(\regs[16][25] ), .B(\regs[17][25] ), .C(\regs[18][25] ), .D(
        \regs[19][25] ), .S0(n1454), .S1(n1430), .Y(n1338) );
  MX4X1 U975 ( .A(\regs[24][25] ), .B(\regs[25][25] ), .C(\regs[26][25] ), .D(
        \regs[27][25] ), .S0(n1454), .S1(n1430), .Y(n1336) );
  MX4X1 U976 ( .A(\regs[20][25] ), .B(\regs[21][25] ), .C(\regs[22][25] ), .D(
        \regs[23][25] ), .S0(n1454), .S1(n1430), .Y(n1337) );
  MX4X1 U977 ( .A(n1388), .B(n1386), .C(n1387), .D(n1385), .S0(n1408), .S1(
        n1410), .Y(n1389) );
  MX4X1 U978 ( .A(\regs[16][30] ), .B(\regs[17][30] ), .C(\regs[18][30] ), .D(
        \regs[19][30] ), .S0(n1457), .S1(n1433), .Y(n1388) );
  MX4X1 U979 ( .A(\regs[24][30] ), .B(\regs[25][30] ), .C(\regs[26][30] ), .D(
        \regs[27][30] ), .S0(n1457), .S1(n1433), .Y(n1386) );
  MX4X1 U980 ( .A(\regs[20][30] ), .B(\regs[21][30] ), .C(\regs[22][30] ), .D(
        \regs[23][30] ), .S0(n1457), .S1(n1433), .Y(n1387) );
  MX4X1 U981 ( .A(n1398), .B(n1396), .C(n1397), .D(n1395), .S0(n1408), .S1(N14), .Y(n1399) );
  MX4X1 U982 ( .A(\regs[16][31] ), .B(\regs[17][31] ), .C(\regs[18][31] ), .D(
        \regs[19][31] ), .S0(n1458), .S1(n1434), .Y(n1398) );
  MX4X1 U983 ( .A(\regs[24][31] ), .B(\regs[25][31] ), .C(\regs[26][31] ), .D(
        \regs[27][31] ), .S0(n1458), .S1(n1434), .Y(n1396) );
  MX4X1 U984 ( .A(\regs[20][31] ), .B(\regs[21][31] ), .C(\regs[22][31] ), .D(
        \regs[23][31] ), .S0(n1458), .S1(n1434), .Y(n1397) );
  MX2X1 U985 ( .A(n1354), .B(n1349), .S0(N16), .Y(N1091) );
  MX4X1 U986 ( .A(n1353), .B(n1351), .C(n1352), .D(n1350), .S0(n1408), .S1(N14), .Y(n1354) );
  MX4X1 U987 ( .A(n1348), .B(n1346), .C(n1347), .D(n1345), .S0(n1408), .S1(N14), .Y(n1349) );
  MX4X1 U988 ( .A(\regs[0][26] ), .B(\regs[1][26] ), .C(\regs[2][26] ), .D(
        \regs[3][26] ), .S0(n1455), .S1(n1431), .Y(n1353) );
  MX2X1 U989 ( .A(n1364), .B(n1359), .S0(N16), .Y(N1090) );
  MX4X1 U990 ( .A(n1363), .B(n1361), .C(n1362), .D(n1360), .S0(n1408), .S1(N14), .Y(n1364) );
  MX4X1 U991 ( .A(n1358), .B(n1356), .C(n1357), .D(n1355), .S0(n1408), .S1(N14), .Y(n1359) );
  MX4X1 U992 ( .A(\regs[0][27] ), .B(\regs[1][27] ), .C(\regs[2][27] ), .D(
        \regs[3][27] ), .S0(n1456), .S1(n1432), .Y(n1363) );
  MX2X1 U993 ( .A(n1374), .B(n1369), .S0(N16), .Y(N1089) );
  MX4X1 U994 ( .A(n1373), .B(n1371), .C(n1372), .D(n1370), .S0(n1408), .S1(
        n1410), .Y(n1374) );
  MX4X1 U995 ( .A(n1368), .B(n1366), .C(n1367), .D(n1365), .S0(n1408), .S1(N14), .Y(n1369) );
  MX4X1 U996 ( .A(\regs[0][28] ), .B(\regs[1][28] ), .C(\regs[2][28] ), .D(
        \regs[3][28] ), .S0(n1456), .S1(n1432), .Y(n1373) );
  MX2X1 U997 ( .A(n1384), .B(n1379), .S0(N16), .Y(N1088) );
  MX4X1 U998 ( .A(n1383), .B(n1381), .C(n1382), .D(n1380), .S0(n1408), .S1(N14), .Y(n1384) );
  MX4X1 U999 ( .A(n1378), .B(n1376), .C(n1377), .D(n1375), .S0(n1408), .S1(N14), .Y(n1379) );
  MX4X1 U1000 ( .A(\regs[0][29] ), .B(\regs[1][29] ), .C(\regs[2][29] ), .D(
        \regs[3][29] ), .S0(n1457), .S1(n1433), .Y(n1383) );
  AND2X2 U1001 ( .A(N1149), .B(reg_ena), .Y(read_data2[0]) );
  MX2X1 U1002 ( .A(n1468), .B(n1463), .S0(N21), .Y(N1149) );
  MX4X1 U1003 ( .A(n1462), .B(n1460), .C(n1461), .D(n1459), .S0(N20), .S1(N19), 
        .Y(n1463) );
  AND2X2 U1004 ( .A(N1148), .B(reg_ena), .Y(read_data2[1]) );
  MX2X1 U1005 ( .A(n1478), .B(n1473), .S0(N21), .Y(N1148) );
  MX4X1 U1006 ( .A(n1477), .B(n1475), .C(n1476), .D(n1474), .S0(N20), .S1(N19), 
        .Y(n1478) );
  AND2X2 U1007 ( .A(N1147), .B(reg_ena), .Y(read_data2[2]) );
  MX2X1 U1008 ( .A(n1488), .B(n1483), .S0(N21), .Y(N1147) );
  MX4X1 U1009 ( .A(n1487), .B(n1485), .C(n1486), .D(n1484), .S0(n1780), .S1(
        n1783), .Y(n1488) );
  AND2X2 U1010 ( .A(N1146), .B(reg_ena), .Y(read_data2[3]) );
  MX2X1 U1011 ( .A(n1498), .B(n1493), .S0(N21), .Y(N1146) );
  MX4X1 U1012 ( .A(n1497), .B(n1495), .C(n1496), .D(n1494), .S0(n1781), .S1(
        n1783), .Y(n1498) );
  AND2X2 U1013 ( .A(N1145), .B(reg_ena), .Y(read_data2[4]) );
  MX2X1 U1014 ( .A(n1508), .B(n1503), .S0(N21), .Y(N1145) );
  MX4X1 U1015 ( .A(n1507), .B(n1505), .C(n1506), .D(n1504), .S0(n1780), .S1(
        n1783), .Y(n1508) );
  AND2X2 U1016 ( .A(N1144), .B(reg_ena), .Y(read_data2[5]) );
  MX2X1 U1017 ( .A(n1518), .B(n1513), .S0(N21), .Y(N1144) );
  MX4X1 U1018 ( .A(n1517), .B(n1515), .C(n1516), .D(n1514), .S0(n1780), .S1(
        n1783), .Y(n1518) );
  AND2X2 U1019 ( .A(N1143), .B(reg_ena), .Y(read_data2[6]) );
  MX2X1 U1020 ( .A(n1528), .B(n1523), .S0(N21), .Y(N1143) );
  MX4X1 U1021 ( .A(n1527), .B(n1525), .C(n1526), .D(n1524), .S0(n1781), .S1(
        n1783), .Y(n1528) );
  AND2X2 U1022 ( .A(N1142), .B(reg_ena), .Y(read_data2[7]) );
  MX2X1 U1023 ( .A(n1538), .B(n1533), .S0(N21), .Y(N1142) );
  MX4X1 U1024 ( .A(n1537), .B(n1535), .C(n1536), .D(n1534), .S0(n1781), .S1(
        n1783), .Y(n1538) );
  AND2X2 U1025 ( .A(N1141), .B(reg_ena), .Y(read_data2[8]) );
  MX2X1 U1026 ( .A(n1548), .B(n1543), .S0(N21), .Y(N1141) );
  MX4X1 U1027 ( .A(n1547), .B(n1545), .C(n1546), .D(n1544), .S0(N20), .S1(
        n1783), .Y(n1548) );
  AND2X2 U1028 ( .A(N1140), .B(reg_ena), .Y(read_data2[9]) );
  MX2X1 U1029 ( .A(n1558), .B(n1553), .S0(N21), .Y(N1140) );
  MX4X1 U1030 ( .A(n1557), .B(n1555), .C(n1556), .D(n1554), .S0(N20), .S1(
        n1783), .Y(n1558) );
  AND2X2 U1031 ( .A(N1139), .B(reg_ena), .Y(read_data2[10]) );
  MX2X1 U1032 ( .A(n1568), .B(n1563), .S0(N21), .Y(N1139) );
  MX4X1 U1033 ( .A(n1567), .B(n1565), .C(n1566), .D(n1564), .S0(n1780), .S1(
        n1783), .Y(n1568) );
  AND2X2 U1034 ( .A(N1138), .B(reg_ena), .Y(read_data2[11]) );
  MX2X1 U1035 ( .A(n1578), .B(n1573), .S0(N21), .Y(N1138) );
  MX4X1 U1036 ( .A(n1577), .B(n1575), .C(n1576), .D(n1574), .S0(N20), .S1(N19), 
        .Y(n1578) );
  AND2X2 U1037 ( .A(N1137), .B(reg_ena), .Y(read_data2[12]) );
  MX2X1 U1038 ( .A(n1588), .B(n1583), .S0(N21), .Y(N1137) );
  MX4X1 U1039 ( .A(n1587), .B(n1585), .C(n1586), .D(n1584), .S0(n1781), .S1(
        n1783), .Y(n1588) );
  AND2X2 U1040 ( .A(N1136), .B(reg_ena), .Y(read_data2[13]) );
  MX2X1 U1041 ( .A(n1598), .B(n1593), .S0(N21), .Y(N1136) );
  MX4X1 U1042 ( .A(n1597), .B(n1595), .C(n1596), .D(n1594), .S0(N20), .S1(N19), 
        .Y(n1598) );
  AND2X2 U1043 ( .A(N1135), .B(reg_ena), .Y(read_data2[14]) );
  MX2X1 U1044 ( .A(n1608), .B(n1603), .S0(N21), .Y(N1135) );
  MX4X1 U1045 ( .A(n1607), .B(n1605), .C(n1606), .D(n1604), .S0(n1780), .S1(
        N19), .Y(n1608) );
  AND2X2 U1046 ( .A(N1134), .B(reg_ena), .Y(read_data2[15]) );
  MX2X1 U1047 ( .A(n1618), .B(n1613), .S0(N21), .Y(N1134) );
  MX4X1 U1048 ( .A(n1617), .B(n1615), .C(n1616), .D(n1614), .S0(n1780), .S1(
        n1783), .Y(n1618) );
  AND2X2 U1049 ( .A(N1133), .B(reg_ena), .Y(read_data2[16]) );
  MX2X1 U1050 ( .A(n1628), .B(n1623), .S0(N21), .Y(N1133) );
  MX4X1 U1051 ( .A(n1627), .B(n1625), .C(n1626), .D(n1624), .S0(n1780), .S1(
        N19), .Y(n1628) );
  AND2X2 U1052 ( .A(N1132), .B(reg_ena), .Y(read_data2[17]) );
  MX2X1 U1053 ( .A(n1638), .B(n1633), .S0(N21), .Y(N1132) );
  MX4X1 U1054 ( .A(n1637), .B(n1635), .C(n1636), .D(n1634), .S0(n1780), .S1(
        N19), .Y(n1638) );
  AND2X2 U1055 ( .A(N1131), .B(reg_ena), .Y(read_data2[18]) );
  MX2X1 U1056 ( .A(n1648), .B(n1643), .S0(N21), .Y(N1131) );
  MX4X1 U1057 ( .A(n1647), .B(n1645), .C(n1646), .D(n1644), .S0(n1780), .S1(
        n1783), .Y(n1648) );
  AND2X2 U1058 ( .A(N1130), .B(reg_ena), .Y(read_data2[19]) );
  MX2X1 U1059 ( .A(n1658), .B(n1653), .S0(N21), .Y(N1130) );
  MX4X1 U1060 ( .A(n1657), .B(n1655), .C(n1656), .D(n1654), .S0(n1780), .S1(
        N19), .Y(n1658) );
  AND2X2 U1061 ( .A(N1129), .B(reg_ena), .Y(read_data2[20]) );
  MX2X1 U1062 ( .A(n1668), .B(n1663), .S0(N21), .Y(N1129) );
  MX4X1 U1063 ( .A(n1667), .B(n1665), .C(n1666), .D(n1664), .S0(n1781), .S1(
        N19), .Y(n1668) );
  AND2X2 U1064 ( .A(N1128), .B(reg_ena), .Y(read_data2[21]) );
  MX2X1 U1065 ( .A(n1678), .B(n1673), .S0(N21), .Y(N1128) );
  MX4X1 U1066 ( .A(n1677), .B(n1675), .C(n1676), .D(n1674), .S0(n1781), .S1(
        N19), .Y(n1678) );
  AND2X2 U1067 ( .A(N1127), .B(reg_ena), .Y(read_data2[22]) );
  MX2X1 U1068 ( .A(n1688), .B(n1683), .S0(N21), .Y(N1127) );
  MX4X1 U1069 ( .A(n1687), .B(n1685), .C(n1686), .D(n1684), .S0(n1781), .S1(
        N19), .Y(n1688) );
  AND2X2 U1070 ( .A(N1126), .B(reg_ena), .Y(read_data2[23]) );
  MX2X1 U1071 ( .A(n1698), .B(n1693), .S0(N21), .Y(N1126) );
  MX4X1 U1072 ( .A(n1697), .B(n1695), .C(n1696), .D(n1694), .S0(n1781), .S1(
        N19), .Y(n1698) );
  AND2X2 U1073 ( .A(N1125), .B(reg_ena), .Y(read_data2[24]) );
  MX2X1 U1074 ( .A(n1708), .B(n1703), .S0(N21), .Y(N1125) );
  MX4X1 U1075 ( .A(n1707), .B(n1705), .C(n1706), .D(n1704), .S0(n1781), .S1(
        N19), .Y(n1708) );
  AND2X2 U1076 ( .A(N1124), .B(reg_ena), .Y(read_data2[25]) );
  MX2X1 U1077 ( .A(n1718), .B(n1713), .S0(N21), .Y(N1124) );
  MX4X1 U1078 ( .A(n1717), .B(n1715), .C(n1716), .D(n1714), .S0(n1781), .S1(
        N19), .Y(n1718) );
  AND2X2 U1079 ( .A(N1123), .B(reg_ena), .Y(read_data2[26]) );
  MX2X1 U1080 ( .A(n1728), .B(n1723), .S0(N21), .Y(N1123) );
  MX4X1 U1081 ( .A(n1727), .B(n1725), .C(n1726), .D(n1724), .S0(N20), .S1(N19), 
        .Y(n1728) );
  AND2X2 U1082 ( .A(N1122), .B(reg_ena), .Y(read_data2[27]) );
  MX2X1 U1083 ( .A(n1738), .B(n1733), .S0(N21), .Y(N1122) );
  MX4X1 U1084 ( .A(n1737), .B(n1735), .C(n1736), .D(n1734), .S0(N20), .S1(N19), 
        .Y(n1738) );
  AND2X2 U1085 ( .A(N1121), .B(reg_ena), .Y(read_data2[28]) );
  MX2X1 U1086 ( .A(n1748), .B(n1743), .S0(N21), .Y(N1121) );
  MX4X1 U1087 ( .A(n1747), .B(n1745), .C(n1746), .D(n1744), .S0(N20), .S1(N19), 
        .Y(n1748) );
  AND2X2 U1088 ( .A(N1120), .B(reg_ena), .Y(read_data2[29]) );
  MX2X1 U1089 ( .A(n1758), .B(n1753), .S0(N21), .Y(N1120) );
  MX4X1 U1090 ( .A(n1757), .B(n1755), .C(n1756), .D(n1754), .S0(N20), .S1(N19), 
        .Y(n1758) );
  AND2X2 U1091 ( .A(N1119), .B(reg_ena), .Y(read_data2[30]) );
  MX2X1 U1092 ( .A(n1768), .B(n1763), .S0(N21), .Y(N1119) );
  MX4X1 U1093 ( .A(n1767), .B(n1765), .C(n1766), .D(n1764), .S0(N20), .S1(N19), 
        .Y(n1768) );
  AND2X2 U1094 ( .A(N1118), .B(reg_ena), .Y(read_data2[31]) );
  MX2X1 U1095 ( .A(n1778), .B(n1773), .S0(N21), .Y(N1118) );
  MX4X1 U1096 ( .A(n1777), .B(n1775), .C(n1776), .D(n1774), .S0(N20), .S1(N19), 
        .Y(n1778) );
  OAI2BB2X1 U1097 ( .B0(n10), .B1(n1), .A0N(\regs[1][7] ), .A1N(n1), .Y(n125)
         );
  OAI2BB2X1 U1098 ( .B0(n11), .B1(n1), .A0N(\regs[1][8] ), .A1N(n1), .Y(n126)
         );
  OAI2BB2X1 U1099 ( .B0(n12), .B1(n1), .A0N(\regs[1][9] ), .A1N(n1), .Y(n127)
         );
  OAI2BB2X1 U1100 ( .B0(n2224), .B1(n1), .A0N(\regs[1][10] ), .A1N(n1), .Y(
        n128) );
  OAI2BB2X1 U1101 ( .B0(n2223), .B1(n1), .A0N(\regs[1][11] ), .A1N(n1), .Y(
        n129) );
  OAI2BB2X1 U1102 ( .B0(n2222), .B1(n1), .A0N(\regs[1][12] ), .A1N(n1), .Y(
        n130) );
  OAI2BB2X1 U1103 ( .B0(n2220), .B1(n1), .A0N(\regs[1][14] ), .A1N(n1), .Y(
        n132) );
  OAI2BB2X1 U1104 ( .B0(n2219), .B1(n1), .A0N(\regs[1][15] ), .A1N(n1), .Y(
        n133) );
  OAI2BB2X1 U1105 ( .B0(n10), .B1(n3), .A0N(\regs[2][7] ), .A1N(n3), .Y(n157)
         );
  OAI2BB2X1 U1106 ( .B0(n11), .B1(n3), .A0N(\regs[2][8] ), .A1N(n3), .Y(n158)
         );
  OAI2BB2X1 U1107 ( .B0(n12), .B1(n3), .A0N(\regs[2][9] ), .A1N(n3), .Y(n159)
         );
  OAI2BB2X1 U1108 ( .B0(n2224), .B1(n3), .A0N(\regs[2][10] ), .A1N(n3), .Y(
        n160) );
  OAI2BB2X1 U1109 ( .B0(n2223), .B1(n3), .A0N(\regs[2][11] ), .A1N(n3), .Y(
        n161) );
  OAI2BB2X1 U1110 ( .B0(n2222), .B1(n3), .A0N(\regs[2][12] ), .A1N(n3), .Y(
        n162) );
  OAI2BB2X1 U1111 ( .B0(n2220), .B1(n3), .A0N(\regs[2][14] ), .A1N(n3), .Y(
        n164) );
  OAI2BB2X1 U1112 ( .B0(n2219), .B1(n3), .A0N(\regs[2][15] ), .A1N(n3), .Y(
        n165) );
  OAI2BB2X1 U1113 ( .B0(n10), .B1(n4), .A0N(\regs[3][7] ), .A1N(n4), .Y(n189)
         );
  OAI2BB2X1 U1114 ( .B0(n11), .B1(n4), .A0N(\regs[3][8] ), .A1N(n4), .Y(n190)
         );
  OAI2BB2X1 U1115 ( .B0(n12), .B1(n4), .A0N(\regs[3][9] ), .A1N(n4), .Y(n191)
         );
  OAI2BB2X1 U1116 ( .B0(n2224), .B1(n4), .A0N(\regs[3][10] ), .A1N(n4), .Y(
        n192) );
  OAI2BB2X1 U1117 ( .B0(n2223), .B1(n4), .A0N(\regs[3][11] ), .A1N(n4), .Y(
        n193) );
  OAI2BB2X1 U1118 ( .B0(n2222), .B1(n4), .A0N(\regs[3][12] ), .A1N(n4), .Y(
        n194) );
  OAI2BB2X1 U1119 ( .B0(n2220), .B1(n4), .A0N(\regs[3][14] ), .A1N(n4), .Y(
        n196) );
  OAI2BB2X1 U1120 ( .B0(n2219), .B1(n4), .A0N(\regs[3][15] ), .A1N(n4), .Y(
        n197) );
  OAI2BB2X1 U1121 ( .B0(n10), .B1(n5), .A0N(\regs[4][7] ), .A1N(n5), .Y(n221)
         );
  OAI2BB2X1 U1122 ( .B0(n11), .B1(n5), .A0N(\regs[4][8] ), .A1N(n5), .Y(n222)
         );
  OAI2BB2X1 U1123 ( .B0(n12), .B1(n5), .A0N(\regs[4][9] ), .A1N(n5), .Y(n223)
         );
  OAI2BB2X1 U1124 ( .B0(n2224), .B1(n5), .A0N(\regs[4][10] ), .A1N(n5), .Y(
        n224) );
  OAI2BB2X1 U1125 ( .B0(n2223), .B1(n5), .A0N(\regs[4][11] ), .A1N(n5), .Y(
        n225) );
  OAI2BB2X1 U1126 ( .B0(n2222), .B1(n5), .A0N(\regs[4][12] ), .A1N(n5), .Y(
        n226) );
  OAI2BB2X1 U1127 ( .B0(n2220), .B1(n5), .A0N(\regs[4][14] ), .A1N(n5), .Y(
        n228) );
  OAI2BB2X1 U1128 ( .B0(n2219), .B1(n5), .A0N(\regs[4][15] ), .A1N(n5), .Y(
        n229) );
  OAI2BB2X1 U1129 ( .B0(n10), .B1(n13), .A0N(\regs[5][7] ), .A1N(n13), .Y(n253) );
  OAI2BB2X1 U1130 ( .B0(n11), .B1(n13), .A0N(\regs[5][8] ), .A1N(n13), .Y(n254) );
  OAI2BB2X1 U1131 ( .B0(n12), .B1(n13), .A0N(\regs[5][9] ), .A1N(n13), .Y(n255) );
  OAI2BB2X1 U1132 ( .B0(n2224), .B1(n13), .A0N(\regs[5][10] ), .A1N(n13), .Y(
        n256) );
  OAI2BB2X1 U1133 ( .B0(n2223), .B1(n13), .A0N(\regs[5][11] ), .A1N(n13), .Y(
        n257) );
  OAI2BB2X1 U1134 ( .B0(n2222), .B1(n13), .A0N(\regs[5][12] ), .A1N(n13), .Y(
        n258) );
  OAI2BB2X1 U1135 ( .B0(n2220), .B1(n13), .A0N(\regs[5][14] ), .A1N(n13), .Y(
        n260) );
  OAI2BB2X1 U1136 ( .B0(n2219), .B1(n13), .A0N(\regs[5][15] ), .A1N(n13), .Y(
        n261) );
  OAI2BB2X1 U1137 ( .B0(n10), .B1(n14), .A0N(\regs[6][7] ), .A1N(n14), .Y(n285) );
  OAI2BB2X1 U1138 ( .B0(n11), .B1(n14), .A0N(\regs[6][8] ), .A1N(n14), .Y(n286) );
  OAI2BB2X1 U1139 ( .B0(n12), .B1(n14), .A0N(\regs[6][9] ), .A1N(n14), .Y(n287) );
  OAI2BB2X1 U1140 ( .B0(n2224), .B1(n14), .A0N(\regs[6][10] ), .A1N(n14), .Y(
        n288) );
  OAI2BB2X1 U1141 ( .B0(n2223), .B1(n14), .A0N(\regs[6][11] ), .A1N(n14), .Y(
        n289) );
  OAI2BB2X1 U1142 ( .B0(n2222), .B1(n14), .A0N(\regs[6][12] ), .A1N(n14), .Y(
        n290) );
  OAI2BB2X1 U1143 ( .B0(n2220), .B1(n14), .A0N(\regs[6][14] ), .A1N(n14), .Y(
        n292) );
  OAI2BB2X1 U1144 ( .B0(n2219), .B1(n14), .A0N(\regs[6][15] ), .A1N(n14), .Y(
        n293) );
  OAI2BB2X1 U1145 ( .B0(n10), .B1(n15), .A0N(\regs[7][7] ), .A1N(n15), .Y(n317) );
  OAI2BB2X1 U1146 ( .B0(n11), .B1(n15), .A0N(\regs[7][8] ), .A1N(n15), .Y(n318) );
  OAI2BB2X1 U1147 ( .B0(n12), .B1(n15), .A0N(\regs[7][9] ), .A1N(n15), .Y(n319) );
  OAI2BB2X1 U1148 ( .B0(n2224), .B1(n15), .A0N(\regs[7][10] ), .A1N(n15), .Y(
        n320) );
  OAI2BB2X1 U1149 ( .B0(n2223), .B1(n15), .A0N(\regs[7][11] ), .A1N(n15), .Y(
        n321) );
  OAI2BB2X1 U1150 ( .B0(n2222), .B1(n15), .A0N(\regs[7][12] ), .A1N(n15), .Y(
        n322) );
  OAI2BB2X1 U1151 ( .B0(n2220), .B1(n15), .A0N(\regs[7][14] ), .A1N(n15), .Y(
        n324) );
  OAI2BB2X1 U1152 ( .B0(n2219), .B1(n15), .A0N(\regs[7][15] ), .A1N(n15), .Y(
        n325) );
  OAI2BB2X1 U1153 ( .B0(n10), .B1(n16), .A0N(\regs[8][7] ), .A1N(n16), .Y(n349) );
  OAI2BB2X1 U1154 ( .B0(n11), .B1(n16), .A0N(\regs[8][8] ), .A1N(n16), .Y(n350) );
  OAI2BB2X1 U1155 ( .B0(n12), .B1(n16), .A0N(\regs[8][9] ), .A1N(n16), .Y(n351) );
  OAI2BB2X1 U1156 ( .B0(n2224), .B1(n16), .A0N(\regs[8][10] ), .A1N(n16), .Y(
        n352) );
  OAI2BB2X1 U1157 ( .B0(n2223), .B1(n16), .A0N(\regs[8][11] ), .A1N(n16), .Y(
        n353) );
  OAI2BB2X1 U1158 ( .B0(n2222), .B1(n16), .A0N(\regs[8][12] ), .A1N(n16), .Y(
        n354) );
  OAI2BB2X1 U1159 ( .B0(n2220), .B1(n16), .A0N(\regs[8][14] ), .A1N(n16), .Y(
        n356) );
  OAI2BB2X1 U1160 ( .B0(n2219), .B1(n16), .A0N(\regs[8][15] ), .A1N(n16), .Y(
        n357) );
  OAI2BB2X1 U1161 ( .B0(n10), .B1(n17), .A0N(\regs[9][7] ), .A1N(n17), .Y(n381) );
  OAI2BB2X1 U1162 ( .B0(n11), .B1(n17), .A0N(\regs[9][8] ), .A1N(n17), .Y(n382) );
  OAI2BB2X1 U1163 ( .B0(n12), .B1(n17), .A0N(\regs[9][9] ), .A1N(n17), .Y(n383) );
  OAI2BB2X1 U1164 ( .B0(n2224), .B1(n17), .A0N(\regs[9][10] ), .A1N(n17), .Y(
        n384) );
  OAI2BB2X1 U1165 ( .B0(n2223), .B1(n17), .A0N(\regs[9][11] ), .A1N(n17), .Y(
        n385) );
  OAI2BB2X1 U1166 ( .B0(n2222), .B1(n17), .A0N(\regs[9][12] ), .A1N(n17), .Y(
        n386) );
  OAI2BB2X1 U1167 ( .B0(n2220), .B1(n17), .A0N(\regs[9][14] ), .A1N(n17), .Y(
        n388) );
  OAI2BB2X1 U1168 ( .B0(n2219), .B1(n17), .A0N(\regs[9][15] ), .A1N(n17), .Y(
        n389) );
  OAI2BB2X1 U1169 ( .B0(n10), .B1(n18), .A0N(\regs[10][7] ), .A1N(n18), .Y(
        n413) );
  OAI2BB2X1 U1170 ( .B0(n11), .B1(n18), .A0N(\regs[10][8] ), .A1N(n18), .Y(
        n414) );
  OAI2BB2X1 U1171 ( .B0(n12), .B1(n18), .A0N(\regs[10][9] ), .A1N(n18), .Y(
        n415) );
  OAI2BB2X1 U1172 ( .B0(n2224), .B1(n18), .A0N(\regs[10][10] ), .A1N(n18), .Y(
        n416) );
  OAI2BB2X1 U1173 ( .B0(n2223), .B1(n18), .A0N(\regs[10][11] ), .A1N(n18), .Y(
        n417) );
  OAI2BB2X1 U1174 ( .B0(n2222), .B1(n18), .A0N(\regs[10][12] ), .A1N(n18), .Y(
        n418) );
  OAI2BB2X1 U1175 ( .B0(n2220), .B1(n18), .A0N(\regs[10][14] ), .A1N(n18), .Y(
        n420) );
  OAI2BB2X1 U1176 ( .B0(n2219), .B1(n18), .A0N(\regs[10][15] ), .A1N(n18), .Y(
        n421) );
  OAI2BB2X1 U1177 ( .B0(n10), .B1(n19), .A0N(\regs[11][7] ), .A1N(n19), .Y(
        n445) );
  OAI2BB2X1 U1178 ( .B0(n11), .B1(n19), .A0N(\regs[11][8] ), .A1N(n19), .Y(
        n446) );
  OAI2BB2X1 U1179 ( .B0(n12), .B1(n19), .A0N(\regs[11][9] ), .A1N(n19), .Y(
        n447) );
  OAI2BB2X1 U1180 ( .B0(n2224), .B1(n19), .A0N(\regs[11][10] ), .A1N(n19), .Y(
        n448) );
  OAI2BB2X1 U1181 ( .B0(n2223), .B1(n19), .A0N(\regs[11][11] ), .A1N(n19), .Y(
        n449) );
  OAI2BB2X1 U1182 ( .B0(n2222), .B1(n19), .A0N(\regs[11][12] ), .A1N(n19), .Y(
        n450) );
  OAI2BB2X1 U1183 ( .B0(n2220), .B1(n19), .A0N(\regs[11][14] ), .A1N(n19), .Y(
        n452) );
  OAI2BB2X1 U1184 ( .B0(n2219), .B1(n19), .A0N(\regs[11][15] ), .A1N(n19), .Y(
        n453) );
  OAI2BB2X1 U1185 ( .B0(n10), .B1(n20), .A0N(\regs[12][7] ), .A1N(n20), .Y(
        n477) );
  OAI2BB2X1 U1186 ( .B0(n11), .B1(n20), .A0N(\regs[12][8] ), .A1N(n20), .Y(
        n478) );
  OAI2BB2X1 U1187 ( .B0(n12), .B1(n20), .A0N(\regs[12][9] ), .A1N(n20), .Y(
        n479) );
  OAI2BB2X1 U1188 ( .B0(n2224), .B1(n20), .A0N(\regs[12][10] ), .A1N(n20), .Y(
        n480) );
  OAI2BB2X1 U1189 ( .B0(n2223), .B1(n20), .A0N(\regs[12][11] ), .A1N(n20), .Y(
        n481) );
  OAI2BB2X1 U1190 ( .B0(n2222), .B1(n20), .A0N(\regs[12][12] ), .A1N(n20), .Y(
        n482) );
  OAI2BB2X1 U1191 ( .B0(n2220), .B1(n20), .A0N(\regs[12][14] ), .A1N(n20), .Y(
        n484) );
  OAI2BB2X1 U1192 ( .B0(n2219), .B1(n20), .A0N(\regs[12][15] ), .A1N(n20), .Y(
        n485) );
  OAI2BB2X1 U1193 ( .B0(n10), .B1(n21), .A0N(\regs[13][7] ), .A1N(n21), .Y(
        n509) );
  OAI2BB2X1 U1194 ( .B0(n11), .B1(n21), .A0N(\regs[13][8] ), .A1N(n21), .Y(
        n510) );
  OAI2BB2X1 U1195 ( .B0(n12), .B1(n21), .A0N(\regs[13][9] ), .A1N(n21), .Y(
        n511) );
  OAI2BB2X1 U1196 ( .B0(n2224), .B1(n21), .A0N(\regs[13][10] ), .A1N(n21), .Y(
        n512) );
  OAI2BB2X1 U1197 ( .B0(n2223), .B1(n21), .A0N(\regs[13][11] ), .A1N(n21), .Y(
        n513) );
  OAI2BB2X1 U1198 ( .B0(n2222), .B1(n21), .A0N(\regs[13][12] ), .A1N(n21), .Y(
        n514) );
  OAI2BB2X1 U1199 ( .B0(n2220), .B1(n21), .A0N(\regs[13][14] ), .A1N(n21), .Y(
        n516) );
  OAI2BB2X1 U1200 ( .B0(n2219), .B1(n21), .A0N(\regs[13][15] ), .A1N(n21), .Y(
        n517) );
  OAI2BB2X1 U1201 ( .B0(n10), .B1(n24), .A0N(\regs[14][7] ), .A1N(n24), .Y(
        n541) );
  OAI2BB2X1 U1202 ( .B0(n11), .B1(n24), .A0N(\regs[14][8] ), .A1N(n24), .Y(
        n542) );
  OAI2BB2X1 U1203 ( .B0(n12), .B1(n24), .A0N(\regs[14][9] ), .A1N(n24), .Y(
        n543) );
  OAI2BB2X1 U1204 ( .B0(n2224), .B1(n24), .A0N(\regs[14][10] ), .A1N(n24), .Y(
        n544) );
  OAI2BB2X1 U1205 ( .B0(n2223), .B1(n24), .A0N(\regs[14][11] ), .A1N(n24), .Y(
        n545) );
  OAI2BB2X1 U1206 ( .B0(n2222), .B1(n24), .A0N(\regs[14][12] ), .A1N(n24), .Y(
        n546) );
  OAI2BB2X1 U1207 ( .B0(n2220), .B1(n24), .A0N(\regs[14][14] ), .A1N(n24), .Y(
        n548) );
  OAI2BB2X1 U1208 ( .B0(n2219), .B1(n24), .A0N(\regs[14][15] ), .A1N(n24), .Y(
        n549) );
  OAI2BB2X1 U1209 ( .B0(n10), .B1(n61), .A0N(\regs[15][7] ), .A1N(n61), .Y(
        n573) );
  OAI2BB2X1 U1210 ( .B0(n11), .B1(n61), .A0N(\regs[15][8] ), .A1N(n61), .Y(
        n574) );
  OAI2BB2X1 U1211 ( .B0(n12), .B1(n61), .A0N(\regs[15][9] ), .A1N(n61), .Y(
        n575) );
  OAI2BB2X1 U1212 ( .B0(n2224), .B1(n61), .A0N(\regs[15][10] ), .A1N(n61), .Y(
        n576) );
  OAI2BB2X1 U1213 ( .B0(n2223), .B1(n61), .A0N(\regs[15][11] ), .A1N(n61), .Y(
        n577) );
  OAI2BB2X1 U1214 ( .B0(n2222), .B1(n61), .A0N(\regs[15][12] ), .A1N(n61), .Y(
        n578) );
  OAI2BB2X1 U1215 ( .B0(n2220), .B1(n61), .A0N(\regs[15][14] ), .A1N(n61), .Y(
        n580) );
  OAI2BB2X1 U1216 ( .B0(n2219), .B1(n61), .A0N(\regs[15][15] ), .A1N(n61), .Y(
        n581) );
  OAI2BB2X1 U1217 ( .B0(n10), .B1(n22), .A0N(\regs[16][7] ), .A1N(n22), .Y(
        n605) );
  OAI2BB2X1 U1218 ( .B0(n11), .B1(n22), .A0N(\regs[16][8] ), .A1N(n22), .Y(
        n606) );
  OAI2BB2X1 U1219 ( .B0(n12), .B1(n22), .A0N(\regs[16][9] ), .A1N(n22), .Y(
        n607) );
  OAI2BB2X1 U1220 ( .B0(n2224), .B1(n22), .A0N(\regs[16][10] ), .A1N(n22), .Y(
        n608) );
  OAI2BB2X1 U1221 ( .B0(n2223), .B1(n22), .A0N(\regs[16][11] ), .A1N(n22), .Y(
        n609) );
  OAI2BB2X1 U1222 ( .B0(n2222), .B1(n22), .A0N(\regs[16][12] ), .A1N(n22), .Y(
        n610) );
  OAI2BB2X1 U1223 ( .B0(n2220), .B1(n22), .A0N(\regs[16][14] ), .A1N(n22), .Y(
        n612) );
  OAI2BB2X1 U1224 ( .B0(n2219), .B1(n22), .A0N(\regs[16][15] ), .A1N(n22), .Y(
        n613) );
  OAI2BB2X1 U1225 ( .B0(n10), .B1(n23), .A0N(\regs[17][7] ), .A1N(n23), .Y(
        n637) );
  OAI2BB2X1 U1226 ( .B0(n11), .B1(n23), .A0N(\regs[17][8] ), .A1N(n23), .Y(
        n638) );
  OAI2BB2X1 U1227 ( .B0(n12), .B1(n23), .A0N(\regs[17][9] ), .A1N(n23), .Y(
        n639) );
  OAI2BB2X1 U1228 ( .B0(n2224), .B1(n23), .A0N(\regs[17][10] ), .A1N(n23), .Y(
        n640) );
  OAI2BB2X1 U1229 ( .B0(n2223), .B1(n23), .A0N(\regs[17][11] ), .A1N(n23), .Y(
        n641) );
  OAI2BB2X1 U1230 ( .B0(n2222), .B1(n23), .A0N(\regs[17][12] ), .A1N(n23), .Y(
        n642) );
  OAI2BB2X1 U1231 ( .B0(n2220), .B1(n23), .A0N(\regs[17][14] ), .A1N(n23), .Y(
        n644) );
  OAI2BB2X1 U1232 ( .B0(n2219), .B1(n23), .A0N(\regs[17][15] ), .A1N(n23), .Y(
        n645) );
  OAI2BB2X1 U1233 ( .B0(n10), .B1(n66), .A0N(\regs[18][7] ), .A1N(n66), .Y(
        n669) );
  OAI2BB2X1 U1234 ( .B0(n11), .B1(n66), .A0N(\regs[18][8] ), .A1N(n66), .Y(
        n670) );
  OAI2BB2X1 U1235 ( .B0(n12), .B1(n66), .A0N(\regs[18][9] ), .A1N(n66), .Y(
        n671) );
  OAI2BB2X1 U1236 ( .B0(n2224), .B1(n66), .A0N(\regs[18][10] ), .A1N(n66), .Y(
        n672) );
  OAI2BB2X1 U1237 ( .B0(n2223), .B1(n66), .A0N(\regs[18][11] ), .A1N(n66), .Y(
        n673) );
  OAI2BB2X1 U1238 ( .B0(n2222), .B1(n66), .A0N(\regs[18][12] ), .A1N(n66), .Y(
        n674) );
  OAI2BB2X1 U1239 ( .B0(n2220), .B1(n66), .A0N(\regs[18][14] ), .A1N(n66), .Y(
        n676) );
  OAI2BB2X1 U1240 ( .B0(n2219), .B1(n66), .A0N(\regs[18][15] ), .A1N(n66), .Y(
        n677) );
  OAI2BB2X1 U1241 ( .B0(n10), .B1(n67), .A0N(\regs[19][7] ), .A1N(n67), .Y(
        n701) );
  OAI2BB2X1 U1242 ( .B0(n11), .B1(n67), .A0N(\regs[19][8] ), .A1N(n67), .Y(
        n702) );
  OAI2BB2X1 U1243 ( .B0(n12), .B1(n67), .A0N(\regs[19][9] ), .A1N(n67), .Y(
        n703) );
  OAI2BB2X1 U1244 ( .B0(n2224), .B1(n67), .A0N(\regs[19][10] ), .A1N(n67), .Y(
        n704) );
  OAI2BB2X1 U1245 ( .B0(n2223), .B1(n67), .A0N(\regs[19][11] ), .A1N(n67), .Y(
        n705) );
  OAI2BB2X1 U1246 ( .B0(n2222), .B1(n67), .A0N(\regs[19][12] ), .A1N(n67), .Y(
        n706) );
  OAI2BB2X1 U1247 ( .B0(n2220), .B1(n67), .A0N(\regs[19][14] ), .A1N(n67), .Y(
        n708) );
  OAI2BB2X1 U1248 ( .B0(n2219), .B1(n67), .A0N(\regs[19][15] ), .A1N(n67), .Y(
        n709) );
  OAI2BB2X1 U1249 ( .B0(n10), .B1(n25), .A0N(\regs[20][7] ), .A1N(n25), .Y(
        n733) );
  OAI2BB2X1 U1250 ( .B0(n11), .B1(n25), .A0N(\regs[20][8] ), .A1N(n25), .Y(
        n734) );
  OAI2BB2X1 U1251 ( .B0(n12), .B1(n25), .A0N(\regs[20][9] ), .A1N(n25), .Y(
        n735) );
  OAI2BB2X1 U1252 ( .B0(n2224), .B1(n25), .A0N(\regs[20][10] ), .A1N(n25), .Y(
        n736) );
  OAI2BB2X1 U1253 ( .B0(n2223), .B1(n25), .A0N(\regs[20][11] ), .A1N(n25), .Y(
        n737) );
  OAI2BB2X1 U1254 ( .B0(n2222), .B1(n25), .A0N(\regs[20][12] ), .A1N(n25), .Y(
        n738) );
  OAI2BB2X1 U1255 ( .B0(n2220), .B1(n25), .A0N(\regs[20][14] ), .A1N(n25), .Y(
        n740) );
  OAI2BB2X1 U1256 ( .B0(n2219), .B1(n25), .A0N(\regs[20][15] ), .A1N(n25), .Y(
        n741) );
  OAI2BB2X1 U1257 ( .B0(n10), .B1(n26), .A0N(\regs[21][7] ), .A1N(n26), .Y(
        n765) );
  OAI2BB2X1 U1258 ( .B0(n11), .B1(n26), .A0N(\regs[21][8] ), .A1N(n26), .Y(
        n766) );
  OAI2BB2X1 U1259 ( .B0(n12), .B1(n26), .A0N(\regs[21][9] ), .A1N(n26), .Y(
        n767) );
  OAI2BB2X1 U1260 ( .B0(n2224), .B1(n26), .A0N(\regs[21][10] ), .A1N(n26), .Y(
        n768) );
  OAI2BB2X1 U1261 ( .B0(n2223), .B1(n26), .A0N(\regs[21][11] ), .A1N(n26), .Y(
        n769) );
  OAI2BB2X1 U1262 ( .B0(n2222), .B1(n26), .A0N(\regs[21][12] ), .A1N(n26), .Y(
        n770) );
  OAI2BB2X1 U1263 ( .B0(n2220), .B1(n26), .A0N(\regs[21][14] ), .A1N(n26), .Y(
        n772) );
  OAI2BB2X1 U1264 ( .B0(n2219), .B1(n26), .A0N(\regs[21][15] ), .A1N(n26), .Y(
        n773) );
  OAI2BB2X1 U1265 ( .B0(n10), .B1(n27), .A0N(\regs[22][7] ), .A1N(n27), .Y(
        n797) );
  OAI2BB2X1 U1266 ( .B0(n11), .B1(n27), .A0N(\regs[22][8] ), .A1N(n27), .Y(
        n798) );
  OAI2BB2X1 U1267 ( .B0(n12), .B1(n27), .A0N(\regs[22][9] ), .A1N(n27), .Y(
        n799) );
  OAI2BB2X1 U1268 ( .B0(n2224), .B1(n27), .A0N(\regs[22][10] ), .A1N(n27), .Y(
        n800) );
  OAI2BB2X1 U1269 ( .B0(n2223), .B1(n27), .A0N(\regs[22][11] ), .A1N(n27), .Y(
        n801) );
  OAI2BB2X1 U1270 ( .B0(n2222), .B1(n27), .A0N(\regs[22][12] ), .A1N(n27), .Y(
        n802) );
  OAI2BB2X1 U1271 ( .B0(n2220), .B1(n27), .A0N(\regs[22][14] ), .A1N(n27), .Y(
        n804) );
  OAI2BB2X1 U1272 ( .B0(n2219), .B1(n27), .A0N(\regs[22][15] ), .A1N(n27), .Y(
        n805) );
  OAI2BB2X1 U1273 ( .B0(n10), .B1(n28), .A0N(\regs[23][7] ), .A1N(n28), .Y(
        n829) );
  OAI2BB2X1 U1274 ( .B0(n11), .B1(n28), .A0N(\regs[23][8] ), .A1N(n28), .Y(
        n830) );
  OAI2BB2X1 U1275 ( .B0(n12), .B1(n28), .A0N(\regs[23][9] ), .A1N(n28), .Y(
        n831) );
  OAI2BB2X1 U1276 ( .B0(n2224), .B1(n28), .A0N(\regs[23][10] ), .A1N(n28), .Y(
        n832) );
  OAI2BB2X1 U1277 ( .B0(n2223), .B1(n28), .A0N(\regs[23][11] ), .A1N(n28), .Y(
        n833) );
  OAI2BB2X1 U1278 ( .B0(n2222), .B1(n28), .A0N(\regs[23][12] ), .A1N(n28), .Y(
        n834) );
  OAI2BB2X1 U1279 ( .B0(n2220), .B1(n28), .A0N(\regs[23][14] ), .A1N(n28), .Y(
        n836) );
  OAI2BB2X1 U1280 ( .B0(n2219), .B1(n28), .A0N(\regs[23][15] ), .A1N(n28), .Y(
        n837) );
  OAI2BB2X1 U1281 ( .B0(n10), .B1(n29), .A0N(\regs[24][7] ), .A1N(n29), .Y(
        n861) );
  OAI2BB2X1 U1282 ( .B0(n11), .B1(n29), .A0N(\regs[24][8] ), .A1N(n29), .Y(
        n862) );
  OAI2BB2X1 U1283 ( .B0(n12), .B1(n29), .A0N(\regs[24][9] ), .A1N(n29), .Y(
        n863) );
  OAI2BB2X1 U1284 ( .B0(n2224), .B1(n29), .A0N(\regs[24][10] ), .A1N(n29), .Y(
        n864) );
  OAI2BB2X1 U1285 ( .B0(n2223), .B1(n29), .A0N(\regs[24][11] ), .A1N(n29), .Y(
        n865) );
  OAI2BB2X1 U1286 ( .B0(n2222), .B1(n29), .A0N(\regs[24][12] ), .A1N(n29), .Y(
        n866) );
  OAI2BB2X1 U1287 ( .B0(n2220), .B1(n29), .A0N(\regs[24][14] ), .A1N(n29), .Y(
        n868) );
  OAI2BB2X1 U1288 ( .B0(n2219), .B1(n29), .A0N(\regs[24][15] ), .A1N(n29), .Y(
        n869) );
  OAI2BB2X1 U1289 ( .B0(n10), .B1(n30), .A0N(\regs[25][7] ), .A1N(n30), .Y(
        n893) );
  OAI2BB2X1 U1290 ( .B0(n11), .B1(n30), .A0N(\regs[25][8] ), .A1N(n30), .Y(
        n894) );
  OAI2BB2X1 U1291 ( .B0(n12), .B1(n30), .A0N(\regs[25][9] ), .A1N(n30), .Y(
        n895) );
  OAI2BB2X1 U1292 ( .B0(n2224), .B1(n30), .A0N(\regs[25][10] ), .A1N(n30), .Y(
        n896) );
  OAI2BB2X1 U1293 ( .B0(n2223), .B1(n30), .A0N(\regs[25][11] ), .A1N(n30), .Y(
        n897) );
  OAI2BB2X1 U1294 ( .B0(n2222), .B1(n30), .A0N(\regs[25][12] ), .A1N(n30), .Y(
        n898) );
  OAI2BB2X1 U1295 ( .B0(n2220), .B1(n30), .A0N(\regs[25][14] ), .A1N(n30), .Y(
        n900) );
  OAI2BB2X1 U1296 ( .B0(n2219), .B1(n30), .A0N(\regs[25][15] ), .A1N(n30), .Y(
        n901) );
  OAI2BB2X1 U1297 ( .B0(n10), .B1(n31), .A0N(\regs[26][7] ), .A1N(n31), .Y(
        n925) );
  OAI2BB2X1 U1298 ( .B0(n11), .B1(n31), .A0N(\regs[26][8] ), .A1N(n31), .Y(
        n926) );
  OAI2BB2X1 U1299 ( .B0(n12), .B1(n31), .A0N(\regs[26][9] ), .A1N(n31), .Y(
        n927) );
  OAI2BB2X1 U1300 ( .B0(n2224), .B1(n31), .A0N(\regs[26][10] ), .A1N(n31), .Y(
        n928) );
  OAI2BB2X1 U1301 ( .B0(n2223), .B1(n31), .A0N(\regs[26][11] ), .A1N(n31), .Y(
        n929) );
  OAI2BB2X1 U1302 ( .B0(n2222), .B1(n31), .A0N(\regs[26][12] ), .A1N(n31), .Y(
        n930) );
  OAI2BB2X1 U1303 ( .B0(n2220), .B1(n31), .A0N(\regs[26][14] ), .A1N(n31), .Y(
        n932) );
  OAI2BB2X1 U1304 ( .B0(n2219), .B1(n31), .A0N(\regs[26][15] ), .A1N(n31), .Y(
        n933) );
  OAI2BB2X1 U1305 ( .B0(n10), .B1(n32), .A0N(\regs[27][7] ), .A1N(n32), .Y(
        n957) );
  OAI2BB2X1 U1306 ( .B0(n11), .B1(n32), .A0N(\regs[27][8] ), .A1N(n32), .Y(
        n958) );
  OAI2BB2X1 U1307 ( .B0(n12), .B1(n32), .A0N(\regs[27][9] ), .A1N(n32), .Y(
        n959) );
  OAI2BB2X1 U1308 ( .B0(n2224), .B1(n32), .A0N(\regs[27][10] ), .A1N(n32), .Y(
        n960) );
  OAI2BB2X1 U1309 ( .B0(n2223), .B1(n32), .A0N(\regs[27][11] ), .A1N(n32), .Y(
        n961) );
  OAI2BB2X1 U1310 ( .B0(n2222), .B1(n32), .A0N(\regs[27][12] ), .A1N(n32), .Y(
        n962) );
  OAI2BB2X1 U1311 ( .B0(n2220), .B1(n32), .A0N(\regs[27][14] ), .A1N(n32), .Y(
        n964) );
  OAI2BB2X1 U1312 ( .B0(n2219), .B1(n32), .A0N(\regs[27][15] ), .A1N(n32), .Y(
        n965) );
  OAI2BB2X1 U1313 ( .B0(n10), .B1(n33), .A0N(\regs[28][7] ), .A1N(n33), .Y(
        n989) );
  OAI2BB2X1 U1314 ( .B0(n11), .B1(n33), .A0N(\regs[28][8] ), .A1N(n33), .Y(
        n990) );
  OAI2BB2X1 U1315 ( .B0(n12), .B1(n33), .A0N(\regs[28][9] ), .A1N(n33), .Y(
        n991) );
  OAI2BB2X1 U1316 ( .B0(n2224), .B1(n33), .A0N(\regs[28][10] ), .A1N(n33), .Y(
        n992) );
  OAI2BB2X1 U1317 ( .B0(n2223), .B1(n33), .A0N(\regs[28][11] ), .A1N(n33), .Y(
        n993) );
  OAI2BB2X1 U1318 ( .B0(n2222), .B1(n33), .A0N(\regs[28][12] ), .A1N(n33), .Y(
        n994) );
  OAI2BB2X1 U1319 ( .B0(n2220), .B1(n33), .A0N(\regs[28][14] ), .A1N(n33), .Y(
        n996) );
  OAI2BB2X1 U1320 ( .B0(n2219), .B1(n33), .A0N(\regs[28][15] ), .A1N(n33), .Y(
        n997) );
  OAI2BB2X1 U1321 ( .B0(n10), .B1(n37), .A0N(\regs[29][7] ), .A1N(n37), .Y(
        n1021) );
  OAI2BB2X1 U1322 ( .B0(n11), .B1(n37), .A0N(\regs[29][8] ), .A1N(n37), .Y(
        n1022) );
  OAI2BB2X1 U1323 ( .B0(n12), .B1(n37), .A0N(\regs[29][9] ), .A1N(n37), .Y(
        n1023) );
  OAI2BB2X1 U1324 ( .B0(n2224), .B1(n37), .A0N(\regs[29][10] ), .A1N(n37), .Y(
        n1024) );
  OAI2BB2X1 U1325 ( .B0(n2223), .B1(n37), .A0N(\regs[29][11] ), .A1N(n37), .Y(
        n1025) );
  OAI2BB2X1 U1326 ( .B0(n2222), .B1(n37), .A0N(\regs[29][12] ), .A1N(n37), .Y(
        n1026) );
  OAI2BB2X1 U1327 ( .B0(n2220), .B1(n37), .A0N(\regs[29][14] ), .A1N(n37), .Y(
        n1028) );
  OAI2BB2X1 U1328 ( .B0(n2219), .B1(n37), .A0N(\regs[29][15] ), .A1N(n37), .Y(
        n1029) );
  OAI2BB2X1 U1329 ( .B0(n10), .B1(n39), .A0N(\regs[30][7] ), .A1N(n39), .Y(
        n1053) );
  OAI2BB2X1 U1330 ( .B0(n11), .B1(n39), .A0N(\regs[30][8] ), .A1N(n39), .Y(
        n1054) );
  OAI2BB2X1 U1331 ( .B0(n12), .B1(n39), .A0N(\regs[30][9] ), .A1N(n39), .Y(
        n1055) );
  OAI2BB2X1 U1332 ( .B0(n2224), .B1(n39), .A0N(\regs[30][10] ), .A1N(n39), .Y(
        n1056) );
  OAI2BB2X1 U1333 ( .B0(n2223), .B1(n39), .A0N(\regs[30][11] ), .A1N(n39), .Y(
        n1057) );
  OAI2BB2X1 U1334 ( .B0(n2222), .B1(n39), .A0N(\regs[30][12] ), .A1N(n39), .Y(
        n1058) );
  OAI2BB2X1 U1335 ( .B0(n2220), .B1(n39), .A0N(\regs[30][14] ), .A1N(n39), .Y(
        n1060) );
  OAI2BB2X1 U1336 ( .B0(n2219), .B1(n39), .A0N(\regs[30][15] ), .A1N(n39), .Y(
        n1061) );
  OAI2BB2X1 U1337 ( .B0(n10), .B1(n41), .A0N(\regs[31][7] ), .A1N(n41), .Y(
        n1085) );
  OAI2BB2X1 U1338 ( .B0(n11), .B1(n41), .A0N(\regs[31][8] ), .A1N(n41), .Y(
        n1086) );
  OAI2BB2X1 U1339 ( .B0(n12), .B1(n41), .A0N(\regs[31][9] ), .A1N(n41), .Y(
        n1087) );
  OAI2BB2X1 U1340 ( .B0(n2224), .B1(n41), .A0N(\regs[31][10] ), .A1N(n41), .Y(
        n1088) );
  OAI2BB2X1 U1341 ( .B0(n2223), .B1(n41), .A0N(\regs[31][11] ), .A1N(n41), .Y(
        n1089) );
  OAI2BB2X1 U1342 ( .B0(n2222), .B1(n41), .A0N(\regs[31][12] ), .A1N(n41), .Y(
        n1090) );
  OAI2BB2X1 U1343 ( .B0(n2220), .B1(n41), .A0N(\regs[31][14] ), .A1N(n41), .Y(
        n1092) );
  OAI2BB2X1 U1344 ( .B0(n2219), .B1(n41), .A0N(\regs[31][15] ), .A1N(n41), .Y(
        n1093) );
  OAI2BB2X1 U1345 ( .B0(n2227), .B1(n1), .A0N(\regs[1][0] ), .A1N(n1), .Y(n118) );
  OAI2BB2X1 U1346 ( .B0(n2226), .B1(n1), .A0N(\regs[1][1] ), .A1N(n1), .Y(n119) );
  OAI2BB2X1 U1347 ( .B0(n2225), .B1(n1), .A0N(\regs[1][2] ), .A1N(n1), .Y(n120) );
  OAI2BB2X1 U1348 ( .B0(n6), .B1(n1), .A0N(\regs[1][3] ), .A1N(n1), .Y(n121)
         );
  OAI2BB2X1 U1349 ( .B0(n7), .B1(n1), .A0N(\regs[1][4] ), .A1N(n1), .Y(n122)
         );
  OAI2BB2X1 U1350 ( .B0(n8), .B1(n1), .A0N(\regs[1][5] ), .A1N(n1), .Y(n123)
         );
  OAI2BB2X1 U1351 ( .B0(n9), .B1(n1), .A0N(\regs[1][6] ), .A1N(n1), .Y(n124)
         );
  OAI2BB2X1 U1352 ( .B0(n2221), .B1(n1), .A0N(\regs[1][13] ), .A1N(n1), .Y(
        n131) );
  OAI2BB2X1 U1353 ( .B0(n2218), .B1(n1), .A0N(\regs[1][16] ), .A1N(n1), .Y(
        n134) );
  OAI2BB2X1 U1354 ( .B0(n2217), .B1(n1), .A0N(\regs[1][17] ), .A1N(n1), .Y(
        n135) );
  OAI2BB2X1 U1355 ( .B0(n2216), .B1(n1), .A0N(\regs[1][18] ), .A1N(n1), .Y(
        n136) );
  OAI2BB2X1 U1356 ( .B0(n2215), .B1(n1), .A0N(\regs[1][19] ), .A1N(n1), .Y(
        n137) );
  OAI2BB2X1 U1357 ( .B0(n2214), .B1(n1), .A0N(\regs[1][20] ), .A1N(n1), .Y(
        n138) );
  OAI2BB2X1 U1358 ( .B0(n2213), .B1(n1), .A0N(\regs[1][21] ), .A1N(n1), .Y(
        n139) );
  OAI2BB2X1 U1359 ( .B0(n2212), .B1(n1), .A0N(\regs[1][22] ), .A1N(n1), .Y(
        n140) );
  OAI2BB2X1 U1360 ( .B0(n2211), .B1(n1), .A0N(\regs[1][23] ), .A1N(n1), .Y(
        n141) );
  OAI2BB2X1 U1361 ( .B0(n2210), .B1(n1), .A0N(\regs[1][24] ), .A1N(n1), .Y(
        n142) );
  OAI2BB2X1 U1362 ( .B0(n2209), .B1(n1), .A0N(\regs[1][25] ), .A1N(n1), .Y(
        n143) );
  OAI2BB2X1 U1363 ( .B0(n2208), .B1(n1), .A0N(\regs[1][26] ), .A1N(n1), .Y(
        n144) );
  OAI2BB2X1 U1364 ( .B0(n2207), .B1(n1), .A0N(\regs[1][27] ), .A1N(n1), .Y(
        n145) );
  OAI2BB2X1 U1365 ( .B0(n2206), .B1(n1), .A0N(\regs[1][28] ), .A1N(n1), .Y(
        n146) );
  OAI2BB2X1 U1366 ( .B0(n2205), .B1(n1), .A0N(\regs[1][29] ), .A1N(n1), .Y(
        n147) );
  OAI2BB2X1 U1367 ( .B0(n2204), .B1(n1), .A0N(\regs[1][30] ), .A1N(n1), .Y(
        n148) );
  OAI2BB2X1 U1368 ( .B0(n34), .B1(n1), .A0N(\regs[1][31] ), .A1N(n1), .Y(n149)
         );
  OAI2BB2X1 U1369 ( .B0(n2227), .B1(n3), .A0N(\regs[2][0] ), .A1N(n3), .Y(n150) );
  OAI2BB2X1 U1370 ( .B0(n2226), .B1(n3), .A0N(\regs[2][1] ), .A1N(n3), .Y(n151) );
  OAI2BB2X1 U1371 ( .B0(n2225), .B1(n3), .A0N(\regs[2][2] ), .A1N(n3), .Y(n152) );
  OAI2BB2X1 U1372 ( .B0(n6), .B1(n3), .A0N(\regs[2][3] ), .A1N(n3), .Y(n153)
         );
  OAI2BB2X1 U1373 ( .B0(n7), .B1(n3), .A0N(\regs[2][4] ), .A1N(n3), .Y(n154)
         );
  OAI2BB2X1 U1374 ( .B0(n8), .B1(n3), .A0N(\regs[2][5] ), .A1N(n3), .Y(n155)
         );
  OAI2BB2X1 U1375 ( .B0(n9), .B1(n3), .A0N(\regs[2][6] ), .A1N(n3), .Y(n156)
         );
  OAI2BB2X1 U1376 ( .B0(n2221), .B1(n3), .A0N(\regs[2][13] ), .A1N(n3), .Y(
        n163) );
  OAI2BB2X1 U1377 ( .B0(n2218), .B1(n3), .A0N(\regs[2][16] ), .A1N(n3), .Y(
        n166) );
  OAI2BB2X1 U1378 ( .B0(n2217), .B1(n3), .A0N(\regs[2][17] ), .A1N(n3), .Y(
        n167) );
  OAI2BB2X1 U1379 ( .B0(n2216), .B1(n3), .A0N(\regs[2][18] ), .A1N(n3), .Y(
        n168) );
  OAI2BB2X1 U1380 ( .B0(n2215), .B1(n3), .A0N(\regs[2][19] ), .A1N(n3), .Y(
        n169) );
  OAI2BB2X1 U1381 ( .B0(n2214), .B1(n3), .A0N(\regs[2][20] ), .A1N(n3), .Y(
        n170) );
  OAI2BB2X1 U1382 ( .B0(n2213), .B1(n3), .A0N(\regs[2][21] ), .A1N(n3), .Y(
        n171) );
  OAI2BB2X1 U1383 ( .B0(n2212), .B1(n3), .A0N(\regs[2][22] ), .A1N(n3), .Y(
        n172) );
  OAI2BB2X1 U1384 ( .B0(n2211), .B1(n3), .A0N(\regs[2][23] ), .A1N(n3), .Y(
        n173) );
  OAI2BB2X1 U1385 ( .B0(n2210), .B1(n3), .A0N(\regs[2][24] ), .A1N(n3), .Y(
        n174) );
  OAI2BB2X1 U1386 ( .B0(n2209), .B1(n3), .A0N(\regs[2][25] ), .A1N(n3), .Y(
        n175) );
  OAI2BB2X1 U1387 ( .B0(n2208), .B1(n3), .A0N(\regs[2][26] ), .A1N(n3), .Y(
        n176) );
  OAI2BB2X1 U1388 ( .B0(n2207), .B1(n3), .A0N(\regs[2][27] ), .A1N(n3), .Y(
        n177) );
  OAI2BB2X1 U1389 ( .B0(n2206), .B1(n3), .A0N(\regs[2][28] ), .A1N(n3), .Y(
        n178) );
  OAI2BB2X1 U1390 ( .B0(n2205), .B1(n3), .A0N(\regs[2][29] ), .A1N(n3), .Y(
        n179) );
  OAI2BB2X1 U1391 ( .B0(n2204), .B1(n3), .A0N(\regs[2][30] ), .A1N(n3), .Y(
        n180) );
  OAI2BB2X1 U1392 ( .B0(n34), .B1(n3), .A0N(\regs[2][31] ), .A1N(n3), .Y(n181)
         );
  OAI2BB2X1 U1393 ( .B0(n2227), .B1(n4), .A0N(\regs[3][0] ), .A1N(n4), .Y(n182) );
  OAI2BB2X1 U1394 ( .B0(n2226), .B1(n4), .A0N(\regs[3][1] ), .A1N(n4), .Y(n183) );
  OAI2BB2X1 U1395 ( .B0(n2225), .B1(n4), .A0N(\regs[3][2] ), .A1N(n4), .Y(n184) );
  OAI2BB2X1 U1396 ( .B0(n6), .B1(n4), .A0N(\regs[3][3] ), .A1N(n4), .Y(n185)
         );
  OAI2BB2X1 U1397 ( .B0(n7), .B1(n4), .A0N(\regs[3][4] ), .A1N(n4), .Y(n186)
         );
  OAI2BB2X1 U1398 ( .B0(n8), .B1(n4), .A0N(\regs[3][5] ), .A1N(n4), .Y(n187)
         );
  OAI2BB2X1 U1399 ( .B0(n9), .B1(n4), .A0N(\regs[3][6] ), .A1N(n4), .Y(n188)
         );
  OAI2BB2X1 U1400 ( .B0(n2221), .B1(n4), .A0N(\regs[3][13] ), .A1N(n4), .Y(
        n195) );
  OAI2BB2X1 U1401 ( .B0(n2218), .B1(n4), .A0N(\regs[3][16] ), .A1N(n4), .Y(
        n198) );
  OAI2BB2X1 U1402 ( .B0(n2217), .B1(n4), .A0N(\regs[3][17] ), .A1N(n4), .Y(
        n199) );
  OAI2BB2X1 U1403 ( .B0(n2216), .B1(n4), .A0N(\regs[3][18] ), .A1N(n4), .Y(
        n200) );
  OAI2BB2X1 U1404 ( .B0(n2215), .B1(n4), .A0N(\regs[3][19] ), .A1N(n4), .Y(
        n201) );
  OAI2BB2X1 U1405 ( .B0(n2214), .B1(n4), .A0N(\regs[3][20] ), .A1N(n4), .Y(
        n202) );
  OAI2BB2X1 U1406 ( .B0(n2213), .B1(n4), .A0N(\regs[3][21] ), .A1N(n4), .Y(
        n203) );
  OAI2BB2X1 U1407 ( .B0(n2212), .B1(n4), .A0N(\regs[3][22] ), .A1N(n4), .Y(
        n204) );
  OAI2BB2X1 U1408 ( .B0(n2211), .B1(n4), .A0N(\regs[3][23] ), .A1N(n4), .Y(
        n205) );
  OAI2BB2X1 U1409 ( .B0(n2210), .B1(n4), .A0N(\regs[3][24] ), .A1N(n4), .Y(
        n206) );
  OAI2BB2X1 U1410 ( .B0(n2209), .B1(n4), .A0N(\regs[3][25] ), .A1N(n4), .Y(
        n207) );
  OAI2BB2X1 U1411 ( .B0(n2208), .B1(n4), .A0N(\regs[3][26] ), .A1N(n4), .Y(
        n208) );
  OAI2BB2X1 U1412 ( .B0(n2207), .B1(n4), .A0N(\regs[3][27] ), .A1N(n4), .Y(
        n209) );
  OAI2BB2X1 U1413 ( .B0(n2206), .B1(n4), .A0N(\regs[3][28] ), .A1N(n4), .Y(
        n210) );
  OAI2BB2X1 U1414 ( .B0(n2205), .B1(n4), .A0N(\regs[3][29] ), .A1N(n4), .Y(
        n211) );
  OAI2BB2X1 U1415 ( .B0(n2204), .B1(n4), .A0N(\regs[3][30] ), .A1N(n4), .Y(
        n212) );
  OAI2BB2X1 U1416 ( .B0(n34), .B1(n4), .A0N(\regs[3][31] ), .A1N(n4), .Y(n213)
         );
  OAI2BB2X1 U1417 ( .B0(n2227), .B1(n5), .A0N(\regs[4][0] ), .A1N(n5), .Y(n214) );
  OAI2BB2X1 U1418 ( .B0(n2226), .B1(n5), .A0N(\regs[4][1] ), .A1N(n5), .Y(n215) );
  OAI2BB2X1 U1419 ( .B0(n2225), .B1(n5), .A0N(\regs[4][2] ), .A1N(n5), .Y(n216) );
  OAI2BB2X1 U1420 ( .B0(n6), .B1(n5), .A0N(\regs[4][3] ), .A1N(n5), .Y(n217)
         );
  OAI2BB2X1 U1421 ( .B0(n7), .B1(n5), .A0N(\regs[4][4] ), .A1N(n5), .Y(n218)
         );
  OAI2BB2X1 U1422 ( .B0(n8), .B1(n5), .A0N(\regs[4][5] ), .A1N(n5), .Y(n219)
         );
  OAI2BB2X1 U1423 ( .B0(n9), .B1(n5), .A0N(\regs[4][6] ), .A1N(n5), .Y(n220)
         );
  OAI2BB2X1 U1424 ( .B0(n2221), .B1(n5), .A0N(\regs[4][13] ), .A1N(n5), .Y(
        n227) );
  OAI2BB2X1 U1425 ( .B0(n2218), .B1(n5), .A0N(\regs[4][16] ), .A1N(n5), .Y(
        n230) );
  OAI2BB2X1 U1426 ( .B0(n2217), .B1(n5), .A0N(\regs[4][17] ), .A1N(n5), .Y(
        n231) );
  OAI2BB2X1 U1427 ( .B0(n2216), .B1(n5), .A0N(\regs[4][18] ), .A1N(n5), .Y(
        n232) );
  OAI2BB2X1 U1428 ( .B0(n2215), .B1(n5), .A0N(\regs[4][19] ), .A1N(n5), .Y(
        n233) );
  OAI2BB2X1 U1429 ( .B0(n2214), .B1(n5), .A0N(\regs[4][20] ), .A1N(n5), .Y(
        n234) );
  OAI2BB2X1 U1430 ( .B0(n2213), .B1(n5), .A0N(\regs[4][21] ), .A1N(n5), .Y(
        n235) );
  OAI2BB2X1 U1431 ( .B0(n2212), .B1(n5), .A0N(\regs[4][22] ), .A1N(n5), .Y(
        n236) );
  OAI2BB2X1 U1432 ( .B0(n2211), .B1(n5), .A0N(\regs[4][23] ), .A1N(n5), .Y(
        n237) );
  OAI2BB2X1 U1433 ( .B0(n2210), .B1(n5), .A0N(\regs[4][24] ), .A1N(n5), .Y(
        n238) );
  OAI2BB2X1 U1434 ( .B0(n2209), .B1(n5), .A0N(\regs[4][25] ), .A1N(n5), .Y(
        n239) );
  OAI2BB2X1 U1435 ( .B0(n2208), .B1(n5), .A0N(\regs[4][26] ), .A1N(n5), .Y(
        n240) );
  OAI2BB2X1 U1436 ( .B0(n2207), .B1(n5), .A0N(\regs[4][27] ), .A1N(n5), .Y(
        n241) );
  OAI2BB2X1 U1437 ( .B0(n2206), .B1(n5), .A0N(\regs[4][28] ), .A1N(n5), .Y(
        n242) );
  OAI2BB2X1 U1438 ( .B0(n2205), .B1(n5), .A0N(\regs[4][29] ), .A1N(n5), .Y(
        n243) );
  OAI2BB2X1 U1439 ( .B0(n2204), .B1(n5), .A0N(\regs[4][30] ), .A1N(n5), .Y(
        n244) );
  OAI2BB2X1 U1440 ( .B0(n34), .B1(n5), .A0N(\regs[4][31] ), .A1N(n5), .Y(n245)
         );
  OAI2BB2X1 U1441 ( .B0(n2227), .B1(n13), .A0N(\regs[5][0] ), .A1N(n13), .Y(
        n246) );
  OAI2BB2X1 U1442 ( .B0(n2226), .B1(n13), .A0N(\regs[5][1] ), .A1N(n13), .Y(
        n247) );
  OAI2BB2X1 U1443 ( .B0(n2225), .B1(n13), .A0N(\regs[5][2] ), .A1N(n13), .Y(
        n248) );
  OAI2BB2X1 U1444 ( .B0(n6), .B1(n13), .A0N(\regs[5][3] ), .A1N(n13), .Y(n249)
         );
  OAI2BB2X1 U1445 ( .B0(n7), .B1(n13), .A0N(\regs[5][4] ), .A1N(n13), .Y(n250)
         );
  OAI2BB2X1 U1446 ( .B0(n8), .B1(n13), .A0N(\regs[5][5] ), .A1N(n13), .Y(n251)
         );
  OAI2BB2X1 U1447 ( .B0(n9), .B1(n13), .A0N(\regs[5][6] ), .A1N(n13), .Y(n252)
         );
  OAI2BB2X1 U1448 ( .B0(n2221), .B1(n13), .A0N(\regs[5][13] ), .A1N(n13), .Y(
        n259) );
  OAI2BB2X1 U1449 ( .B0(n2218), .B1(n13), .A0N(\regs[5][16] ), .A1N(n13), .Y(
        n262) );
  OAI2BB2X1 U1450 ( .B0(n2217), .B1(n13), .A0N(\regs[5][17] ), .A1N(n13), .Y(
        n263) );
  OAI2BB2X1 U1451 ( .B0(n2216), .B1(n13), .A0N(\regs[5][18] ), .A1N(n13), .Y(
        n264) );
  OAI2BB2X1 U1452 ( .B0(n2215), .B1(n13), .A0N(\regs[5][19] ), .A1N(n13), .Y(
        n265) );
  OAI2BB2X1 U1453 ( .B0(n2214), .B1(n13), .A0N(\regs[5][20] ), .A1N(n13), .Y(
        n266) );
  OAI2BB2X1 U1454 ( .B0(n2213), .B1(n13), .A0N(\regs[5][21] ), .A1N(n13), .Y(
        n267) );
  OAI2BB2X1 U1455 ( .B0(n2212), .B1(n13), .A0N(\regs[5][22] ), .A1N(n13), .Y(
        n268) );
  OAI2BB2X1 U1456 ( .B0(n2211), .B1(n13), .A0N(\regs[5][23] ), .A1N(n13), .Y(
        n269) );
  OAI2BB2X1 U1457 ( .B0(n2210), .B1(n13), .A0N(\regs[5][24] ), .A1N(n13), .Y(
        n270) );
  OAI2BB2X1 U1458 ( .B0(n2209), .B1(n13), .A0N(\regs[5][25] ), .A1N(n13), .Y(
        n271) );
  OAI2BB2X1 U1459 ( .B0(n2208), .B1(n13), .A0N(\regs[5][26] ), .A1N(n13), .Y(
        n272) );
  OAI2BB2X1 U1460 ( .B0(n2207), .B1(n13), .A0N(\regs[5][27] ), .A1N(n13), .Y(
        n273) );
  OAI2BB2X1 U1461 ( .B0(n2206), .B1(n13), .A0N(\regs[5][28] ), .A1N(n13), .Y(
        n274) );
  OAI2BB2X1 U1462 ( .B0(n2205), .B1(n13), .A0N(\regs[5][29] ), .A1N(n13), .Y(
        n275) );
  OAI2BB2X1 U1463 ( .B0(n2204), .B1(n13), .A0N(\regs[5][30] ), .A1N(n13), .Y(
        n276) );
  OAI2BB2X1 U1464 ( .B0(n34), .B1(n13), .A0N(\regs[5][31] ), .A1N(n13), .Y(
        n277) );
  OAI2BB2X1 U1465 ( .B0(n2227), .B1(n14), .A0N(\regs[6][0] ), .A1N(n14), .Y(
        n278) );
  OAI2BB2X1 U1466 ( .B0(n2226), .B1(n14), .A0N(\regs[6][1] ), .A1N(n14), .Y(
        n279) );
  OAI2BB2X1 U1467 ( .B0(n2225), .B1(n14), .A0N(\regs[6][2] ), .A1N(n14), .Y(
        n280) );
  OAI2BB2X1 U1468 ( .B0(n6), .B1(n14), .A0N(\regs[6][3] ), .A1N(n14), .Y(n281)
         );
  OAI2BB2X1 U1469 ( .B0(n7), .B1(n14), .A0N(\regs[6][4] ), .A1N(n14), .Y(n282)
         );
  OAI2BB2X1 U1470 ( .B0(n8), .B1(n14), .A0N(\regs[6][5] ), .A1N(n14), .Y(n283)
         );
  OAI2BB2X1 U1471 ( .B0(n9), .B1(n14), .A0N(\regs[6][6] ), .A1N(n14), .Y(n284)
         );
  OAI2BB2X1 U1472 ( .B0(n2221), .B1(n14), .A0N(\regs[6][13] ), .A1N(n14), .Y(
        n291) );
  OAI2BB2X1 U1473 ( .B0(n2218), .B1(n14), .A0N(\regs[6][16] ), .A1N(n14), .Y(
        n294) );
  OAI2BB2X1 U1474 ( .B0(n2217), .B1(n14), .A0N(\regs[6][17] ), .A1N(n14), .Y(
        n295) );
  OAI2BB2X1 U1475 ( .B0(n2216), .B1(n14), .A0N(\regs[6][18] ), .A1N(n14), .Y(
        n296) );
  OAI2BB2X1 U1476 ( .B0(n2215), .B1(n14), .A0N(\regs[6][19] ), .A1N(n14), .Y(
        n297) );
  OAI2BB2X1 U1477 ( .B0(n2214), .B1(n14), .A0N(\regs[6][20] ), .A1N(n14), .Y(
        n298) );
  OAI2BB2X1 U1478 ( .B0(n2213), .B1(n14), .A0N(\regs[6][21] ), .A1N(n14), .Y(
        n299) );
  OAI2BB2X1 U1479 ( .B0(n2212), .B1(n14), .A0N(\regs[6][22] ), .A1N(n14), .Y(
        n300) );
  OAI2BB2X1 U1480 ( .B0(n2211), .B1(n14), .A0N(\regs[6][23] ), .A1N(n14), .Y(
        n301) );
  OAI2BB2X1 U1481 ( .B0(n2210), .B1(n14), .A0N(\regs[6][24] ), .A1N(n14), .Y(
        n302) );
  OAI2BB2X1 U1482 ( .B0(n2209), .B1(n14), .A0N(\regs[6][25] ), .A1N(n14), .Y(
        n303) );
  OAI2BB2X1 U1483 ( .B0(n2208), .B1(n14), .A0N(\regs[6][26] ), .A1N(n14), .Y(
        n304) );
  OAI2BB2X1 U1484 ( .B0(n2207), .B1(n14), .A0N(\regs[6][27] ), .A1N(n14), .Y(
        n305) );
  OAI2BB2X1 U1485 ( .B0(n2206), .B1(n14), .A0N(\regs[6][28] ), .A1N(n14), .Y(
        n306) );
  OAI2BB2X1 U1486 ( .B0(n2205), .B1(n14), .A0N(\regs[6][29] ), .A1N(n14), .Y(
        n307) );
  OAI2BB2X1 U1487 ( .B0(n2204), .B1(n14), .A0N(\regs[6][30] ), .A1N(n14), .Y(
        n308) );
  OAI2BB2X1 U1488 ( .B0(n34), .B1(n14), .A0N(\regs[6][31] ), .A1N(n14), .Y(
        n309) );
  OAI2BB2X1 U1489 ( .B0(n2227), .B1(n15), .A0N(\regs[7][0] ), .A1N(n15), .Y(
        n310) );
  OAI2BB2X1 U1490 ( .B0(n2226), .B1(n15), .A0N(\regs[7][1] ), .A1N(n15), .Y(
        n311) );
  OAI2BB2X1 U1491 ( .B0(n2225), .B1(n15), .A0N(\regs[7][2] ), .A1N(n15), .Y(
        n312) );
  OAI2BB2X1 U1492 ( .B0(n6), .B1(n15), .A0N(\regs[7][3] ), .A1N(n15), .Y(n313)
         );
  OAI2BB2X1 U1493 ( .B0(n7), .B1(n15), .A0N(\regs[7][4] ), .A1N(n15), .Y(n314)
         );
  OAI2BB2X1 U1494 ( .B0(n8), .B1(n15), .A0N(\regs[7][5] ), .A1N(n15), .Y(n315)
         );
  OAI2BB2X1 U1495 ( .B0(n9), .B1(n15), .A0N(\regs[7][6] ), .A1N(n15), .Y(n316)
         );
  OAI2BB2X1 U1496 ( .B0(n2221), .B1(n15), .A0N(\regs[7][13] ), .A1N(n15), .Y(
        n323) );
  OAI2BB2X1 U1497 ( .B0(n2218), .B1(n15), .A0N(\regs[7][16] ), .A1N(n15), .Y(
        n326) );
  OAI2BB2X1 U1498 ( .B0(n2217), .B1(n15), .A0N(\regs[7][17] ), .A1N(n15), .Y(
        n327) );
  OAI2BB2X1 U1499 ( .B0(n2216), .B1(n15), .A0N(\regs[7][18] ), .A1N(n15), .Y(
        n328) );
  OAI2BB2X1 U1500 ( .B0(n2215), .B1(n15), .A0N(\regs[7][19] ), .A1N(n15), .Y(
        n329) );
  OAI2BB2X1 U1501 ( .B0(n2214), .B1(n15), .A0N(\regs[7][20] ), .A1N(n15), .Y(
        n330) );
  OAI2BB2X1 U1502 ( .B0(n2213), .B1(n15), .A0N(\regs[7][21] ), .A1N(n15), .Y(
        n331) );
  OAI2BB2X1 U1503 ( .B0(n2212), .B1(n15), .A0N(\regs[7][22] ), .A1N(n15), .Y(
        n332) );
  OAI2BB2X1 U1504 ( .B0(n2211), .B1(n15), .A0N(\regs[7][23] ), .A1N(n15), .Y(
        n333) );
  OAI2BB2X1 U1505 ( .B0(n2210), .B1(n15), .A0N(\regs[7][24] ), .A1N(n15), .Y(
        n334) );
  OAI2BB2X1 U1506 ( .B0(n2209), .B1(n15), .A0N(\regs[7][25] ), .A1N(n15), .Y(
        n335) );
  OAI2BB2X1 U1507 ( .B0(n2208), .B1(n15), .A0N(\regs[7][26] ), .A1N(n15), .Y(
        n336) );
  OAI2BB2X1 U1508 ( .B0(n2207), .B1(n15), .A0N(\regs[7][27] ), .A1N(n15), .Y(
        n337) );
  OAI2BB2X1 U1509 ( .B0(n2206), .B1(n15), .A0N(\regs[7][28] ), .A1N(n15), .Y(
        n338) );
  OAI2BB2X1 U1510 ( .B0(n2205), .B1(n15), .A0N(\regs[7][29] ), .A1N(n15), .Y(
        n339) );
  OAI2BB2X1 U1511 ( .B0(n2204), .B1(n15), .A0N(\regs[7][30] ), .A1N(n15), .Y(
        n340) );
  OAI2BB2X1 U1512 ( .B0(n34), .B1(n15), .A0N(\regs[7][31] ), .A1N(n15), .Y(
        n341) );
  OAI2BB2X1 U1513 ( .B0(n2227), .B1(n16), .A0N(\regs[8][0] ), .A1N(n16), .Y(
        n342) );
  OAI2BB2X1 U1514 ( .B0(n2226), .B1(n16), .A0N(\regs[8][1] ), .A1N(n16), .Y(
        n343) );
  OAI2BB2X1 U1515 ( .B0(n2225), .B1(n16), .A0N(\regs[8][2] ), .A1N(n16), .Y(
        n344) );
  OAI2BB2X1 U1516 ( .B0(n6), .B1(n16), .A0N(\regs[8][3] ), .A1N(n16), .Y(n345)
         );
  OAI2BB2X1 U1517 ( .B0(n7), .B1(n16), .A0N(\regs[8][4] ), .A1N(n16), .Y(n346)
         );
  OAI2BB2X1 U1518 ( .B0(n8), .B1(n16), .A0N(\regs[8][5] ), .A1N(n16), .Y(n347)
         );
  OAI2BB2X1 U1519 ( .B0(n9), .B1(n16), .A0N(\regs[8][6] ), .A1N(n16), .Y(n348)
         );
  OAI2BB2X1 U1520 ( .B0(n2221), .B1(n16), .A0N(\regs[8][13] ), .A1N(n16), .Y(
        n355) );
  OAI2BB2X1 U1521 ( .B0(n2218), .B1(n16), .A0N(\regs[8][16] ), .A1N(n16), .Y(
        n358) );
  OAI2BB2X1 U1522 ( .B0(n2217), .B1(n16), .A0N(\regs[8][17] ), .A1N(n16), .Y(
        n359) );
  OAI2BB2X1 U1523 ( .B0(n2216), .B1(n16), .A0N(\regs[8][18] ), .A1N(n16), .Y(
        n360) );
  OAI2BB2X1 U1524 ( .B0(n2215), .B1(n16), .A0N(\regs[8][19] ), .A1N(n16), .Y(
        n361) );
  OAI2BB2X1 U1525 ( .B0(n2214), .B1(n16), .A0N(\regs[8][20] ), .A1N(n16), .Y(
        n362) );
  OAI2BB2X1 U1526 ( .B0(n2213), .B1(n16), .A0N(\regs[8][21] ), .A1N(n16), .Y(
        n363) );
  OAI2BB2X1 U1527 ( .B0(n2212), .B1(n16), .A0N(\regs[8][22] ), .A1N(n16), .Y(
        n364) );
  OAI2BB2X1 U1528 ( .B0(n2211), .B1(n16), .A0N(\regs[8][23] ), .A1N(n16), .Y(
        n365) );
  OAI2BB2X1 U1529 ( .B0(n2210), .B1(n16), .A0N(\regs[8][24] ), .A1N(n16), .Y(
        n366) );
  OAI2BB2X1 U1530 ( .B0(n2209), .B1(n16), .A0N(\regs[8][25] ), .A1N(n16), .Y(
        n367) );
  OAI2BB2X1 U1531 ( .B0(n2208), .B1(n16), .A0N(\regs[8][26] ), .A1N(n16), .Y(
        n368) );
  OAI2BB2X1 U1532 ( .B0(n2207), .B1(n16), .A0N(\regs[8][27] ), .A1N(n16), .Y(
        n369) );
  OAI2BB2X1 U1533 ( .B0(n2206), .B1(n16), .A0N(\regs[8][28] ), .A1N(n16), .Y(
        n370) );
  OAI2BB2X1 U1534 ( .B0(n2205), .B1(n16), .A0N(\regs[8][29] ), .A1N(n16), .Y(
        n371) );
  OAI2BB2X1 U1535 ( .B0(n2204), .B1(n16), .A0N(\regs[8][30] ), .A1N(n16), .Y(
        n372) );
  OAI2BB2X1 U1536 ( .B0(n34), .B1(n16), .A0N(\regs[8][31] ), .A1N(n16), .Y(
        n373) );
  OAI2BB2X1 U1537 ( .B0(n2227), .B1(n17), .A0N(\regs[9][0] ), .A1N(n17), .Y(
        n374) );
  OAI2BB2X1 U1538 ( .B0(n2226), .B1(n17), .A0N(\regs[9][1] ), .A1N(n17), .Y(
        n375) );
  OAI2BB2X1 U1539 ( .B0(n2225), .B1(n17), .A0N(\regs[9][2] ), .A1N(n17), .Y(
        n376) );
  OAI2BB2X1 U1540 ( .B0(n6), .B1(n17), .A0N(\regs[9][3] ), .A1N(n17), .Y(n377)
         );
  OAI2BB2X1 U1541 ( .B0(n7), .B1(n17), .A0N(\regs[9][4] ), .A1N(n17), .Y(n378)
         );
  OAI2BB2X1 U1542 ( .B0(n8), .B1(n17), .A0N(\regs[9][5] ), .A1N(n17), .Y(n379)
         );
  OAI2BB2X1 U1543 ( .B0(n9), .B1(n17), .A0N(\regs[9][6] ), .A1N(n17), .Y(n380)
         );
  OAI2BB2X1 U1544 ( .B0(n2221), .B1(n17), .A0N(\regs[9][13] ), .A1N(n17), .Y(
        n387) );
  OAI2BB2X1 U1545 ( .B0(n2218), .B1(n17), .A0N(\regs[9][16] ), .A1N(n17), .Y(
        n390) );
  OAI2BB2X1 U1546 ( .B0(n2217), .B1(n17), .A0N(\regs[9][17] ), .A1N(n17), .Y(
        n391) );
  OAI2BB2X1 U1547 ( .B0(n2216), .B1(n17), .A0N(\regs[9][18] ), .A1N(n17), .Y(
        n392) );
  OAI2BB2X1 U1548 ( .B0(n2215), .B1(n17), .A0N(\regs[9][19] ), .A1N(n17), .Y(
        n393) );
  OAI2BB2X1 U1549 ( .B0(n2214), .B1(n17), .A0N(\regs[9][20] ), .A1N(n17), .Y(
        n394) );
  OAI2BB2X1 U1550 ( .B0(n2213), .B1(n17), .A0N(\regs[9][21] ), .A1N(n17), .Y(
        n395) );
  OAI2BB2X1 U1551 ( .B0(n2212), .B1(n17), .A0N(\regs[9][22] ), .A1N(n17), .Y(
        n396) );
  OAI2BB2X1 U1552 ( .B0(n2211), .B1(n17), .A0N(\regs[9][23] ), .A1N(n17), .Y(
        n397) );
  OAI2BB2X1 U1553 ( .B0(n2210), .B1(n17), .A0N(\regs[9][24] ), .A1N(n17), .Y(
        n398) );
  OAI2BB2X1 U1554 ( .B0(n2209), .B1(n17), .A0N(\regs[9][25] ), .A1N(n17), .Y(
        n399) );
  OAI2BB2X1 U1555 ( .B0(n2208), .B1(n17), .A0N(\regs[9][26] ), .A1N(n17), .Y(
        n400) );
  OAI2BB2X1 U1556 ( .B0(n2207), .B1(n17), .A0N(\regs[9][27] ), .A1N(n17), .Y(
        n401) );
  OAI2BB2X1 U1557 ( .B0(n2206), .B1(n17), .A0N(\regs[9][28] ), .A1N(n17), .Y(
        n402) );
  OAI2BB2X1 U1558 ( .B0(n2205), .B1(n17), .A0N(\regs[9][29] ), .A1N(n17), .Y(
        n403) );
  OAI2BB2X1 U1559 ( .B0(n2204), .B1(n17), .A0N(\regs[9][30] ), .A1N(n17), .Y(
        n404) );
  OAI2BB2X1 U1560 ( .B0(n34), .B1(n17), .A0N(\regs[9][31] ), .A1N(n17), .Y(
        n405) );
  OAI2BB2X1 U1561 ( .B0(n2227), .B1(n18), .A0N(\regs[10][0] ), .A1N(n18), .Y(
        n406) );
  OAI2BB2X1 U1562 ( .B0(n2226), .B1(n18), .A0N(\regs[10][1] ), .A1N(n18), .Y(
        n407) );
  OAI2BB2X1 U1563 ( .B0(n2225), .B1(n18), .A0N(\regs[10][2] ), .A1N(n18), .Y(
        n408) );
  OAI2BB2X1 U1564 ( .B0(n6), .B1(n18), .A0N(\regs[10][3] ), .A1N(n18), .Y(n409) );
  OAI2BB2X1 U1565 ( .B0(n7), .B1(n18), .A0N(\regs[10][4] ), .A1N(n18), .Y(n410) );
  OAI2BB2X1 U1566 ( .B0(n8), .B1(n18), .A0N(\regs[10][5] ), .A1N(n18), .Y(n411) );
  OAI2BB2X1 U1567 ( .B0(n9), .B1(n18), .A0N(\regs[10][6] ), .A1N(n18), .Y(n412) );
  OAI2BB2X1 U1568 ( .B0(n2221), .B1(n18), .A0N(\regs[10][13] ), .A1N(n18), .Y(
        n419) );
  OAI2BB2X1 U1569 ( .B0(n2218), .B1(n18), .A0N(\regs[10][16] ), .A1N(n18), .Y(
        n422) );
  OAI2BB2X1 U1570 ( .B0(n2217), .B1(n18), .A0N(\regs[10][17] ), .A1N(n18), .Y(
        n423) );
  OAI2BB2X1 U1571 ( .B0(n2216), .B1(n18), .A0N(\regs[10][18] ), .A1N(n18), .Y(
        n424) );
  OAI2BB2X1 U1572 ( .B0(n2215), .B1(n18), .A0N(\regs[10][19] ), .A1N(n18), .Y(
        n425) );
  OAI2BB2X1 U1573 ( .B0(n2214), .B1(n18), .A0N(\regs[10][20] ), .A1N(n18), .Y(
        n426) );
  OAI2BB2X1 U1574 ( .B0(n2213), .B1(n18), .A0N(\regs[10][21] ), .A1N(n18), .Y(
        n427) );
  OAI2BB2X1 U1575 ( .B0(n2212), .B1(n18), .A0N(\regs[10][22] ), .A1N(n18), .Y(
        n428) );
  OAI2BB2X1 U1576 ( .B0(n2211), .B1(n18), .A0N(\regs[10][23] ), .A1N(n18), .Y(
        n429) );
  OAI2BB2X1 U1577 ( .B0(n2210), .B1(n18), .A0N(\regs[10][24] ), .A1N(n18), .Y(
        n430) );
  OAI2BB2X1 U1578 ( .B0(n2209), .B1(n18), .A0N(\regs[10][25] ), .A1N(n18), .Y(
        n431) );
  OAI2BB2X1 U1579 ( .B0(n2208), .B1(n18), .A0N(\regs[10][26] ), .A1N(n18), .Y(
        n432) );
  OAI2BB2X1 U1580 ( .B0(n2207), .B1(n18), .A0N(\regs[10][27] ), .A1N(n18), .Y(
        n433) );
  OAI2BB2X1 U1581 ( .B0(n2206), .B1(n18), .A0N(\regs[10][28] ), .A1N(n18), .Y(
        n434) );
  OAI2BB2X1 U1582 ( .B0(n2205), .B1(n18), .A0N(\regs[10][29] ), .A1N(n18), .Y(
        n435) );
  OAI2BB2X1 U1583 ( .B0(n2204), .B1(n18), .A0N(\regs[10][30] ), .A1N(n18), .Y(
        n436) );
  OAI2BB2X1 U1584 ( .B0(n34), .B1(n18), .A0N(\regs[10][31] ), .A1N(n18), .Y(
        n437) );
  OAI2BB2X1 U1585 ( .B0(n2227), .B1(n19), .A0N(\regs[11][0] ), .A1N(n19), .Y(
        n438) );
  OAI2BB2X1 U1586 ( .B0(n2226), .B1(n19), .A0N(\regs[11][1] ), .A1N(n19), .Y(
        n439) );
  OAI2BB2X1 U1587 ( .B0(n2225), .B1(n19), .A0N(\regs[11][2] ), .A1N(n19), .Y(
        n440) );
  OAI2BB2X1 U1588 ( .B0(n6), .B1(n19), .A0N(\regs[11][3] ), .A1N(n19), .Y(n441) );
  OAI2BB2X1 U1589 ( .B0(n7), .B1(n19), .A0N(\regs[11][4] ), .A1N(n19), .Y(n442) );
  OAI2BB2X1 U1590 ( .B0(n8), .B1(n19), .A0N(\regs[11][5] ), .A1N(n19), .Y(n443) );
  OAI2BB2X1 U1591 ( .B0(n9), .B1(n19), .A0N(\regs[11][6] ), .A1N(n19), .Y(n444) );
  OAI2BB2X1 U1592 ( .B0(n2221), .B1(n19), .A0N(\regs[11][13] ), .A1N(n19), .Y(
        n451) );
  OAI2BB2X1 U1593 ( .B0(n2218), .B1(n19), .A0N(\regs[11][16] ), .A1N(n19), .Y(
        n454) );
  OAI2BB2X1 U1594 ( .B0(n2217), .B1(n19), .A0N(\regs[11][17] ), .A1N(n19), .Y(
        n455) );
  OAI2BB2X1 U1595 ( .B0(n2216), .B1(n19), .A0N(\regs[11][18] ), .A1N(n19), .Y(
        n456) );
  OAI2BB2X1 U1596 ( .B0(n2215), .B1(n19), .A0N(\regs[11][19] ), .A1N(n19), .Y(
        n457) );
  OAI2BB2X1 U1597 ( .B0(n2214), .B1(n19), .A0N(\regs[11][20] ), .A1N(n19), .Y(
        n458) );
  OAI2BB2X1 U1598 ( .B0(n2213), .B1(n19), .A0N(\regs[11][21] ), .A1N(n19), .Y(
        n459) );
  OAI2BB2X1 U1599 ( .B0(n2212), .B1(n19), .A0N(\regs[11][22] ), .A1N(n19), .Y(
        n460) );
  OAI2BB2X1 U1600 ( .B0(n2211), .B1(n19), .A0N(\regs[11][23] ), .A1N(n19), .Y(
        n461) );
  OAI2BB2X1 U1601 ( .B0(n2210), .B1(n19), .A0N(\regs[11][24] ), .A1N(n19), .Y(
        n462) );
  OAI2BB2X1 U1602 ( .B0(n2209), .B1(n19), .A0N(\regs[11][25] ), .A1N(n19), .Y(
        n463) );
  OAI2BB2X1 U1603 ( .B0(n2208), .B1(n19), .A0N(\regs[11][26] ), .A1N(n19), .Y(
        n464) );
  OAI2BB2X1 U1604 ( .B0(n2207), .B1(n19), .A0N(\regs[11][27] ), .A1N(n19), .Y(
        n465) );
  OAI2BB2X1 U1605 ( .B0(n2206), .B1(n19), .A0N(\regs[11][28] ), .A1N(n19), .Y(
        n466) );
  OAI2BB2X1 U1606 ( .B0(n2205), .B1(n19), .A0N(\regs[11][29] ), .A1N(n19), .Y(
        n467) );
  OAI2BB2X1 U1607 ( .B0(n2204), .B1(n19), .A0N(\regs[11][30] ), .A1N(n19), .Y(
        n468) );
  OAI2BB2X1 U1608 ( .B0(n34), .B1(n19), .A0N(\regs[11][31] ), .A1N(n19), .Y(
        n469) );
  OAI2BB2X1 U1609 ( .B0(n2227), .B1(n20), .A0N(\regs[12][0] ), .A1N(n20), .Y(
        n470) );
  OAI2BB2X1 U1610 ( .B0(n2226), .B1(n20), .A0N(\regs[12][1] ), .A1N(n20), .Y(
        n471) );
  OAI2BB2X1 U1611 ( .B0(n2225), .B1(n20), .A0N(\regs[12][2] ), .A1N(n20), .Y(
        n472) );
  OAI2BB2X1 U1612 ( .B0(n6), .B1(n20), .A0N(\regs[12][3] ), .A1N(n20), .Y(n473) );
  OAI2BB2X1 U1613 ( .B0(n7), .B1(n20), .A0N(\regs[12][4] ), .A1N(n20), .Y(n474) );
  OAI2BB2X1 U1614 ( .B0(n8), .B1(n20), .A0N(\regs[12][5] ), .A1N(n20), .Y(n475) );
  OAI2BB2X1 U1615 ( .B0(n9), .B1(n20), .A0N(\regs[12][6] ), .A1N(n20), .Y(n476) );
  OAI2BB2X1 U1616 ( .B0(n2221), .B1(n20), .A0N(\regs[12][13] ), .A1N(n20), .Y(
        n483) );
  OAI2BB2X1 U1617 ( .B0(n2218), .B1(n20), .A0N(\regs[12][16] ), .A1N(n20), .Y(
        n486) );
  OAI2BB2X1 U1618 ( .B0(n2217), .B1(n20), .A0N(\regs[12][17] ), .A1N(n20), .Y(
        n487) );
  OAI2BB2X1 U1619 ( .B0(n2216), .B1(n20), .A0N(\regs[12][18] ), .A1N(n20), .Y(
        n488) );
  OAI2BB2X1 U1620 ( .B0(n2215), .B1(n20), .A0N(\regs[12][19] ), .A1N(n20), .Y(
        n489) );
  OAI2BB2X1 U1621 ( .B0(n2214), .B1(n20), .A0N(\regs[12][20] ), .A1N(n20), .Y(
        n490) );
  OAI2BB2X1 U1622 ( .B0(n2213), .B1(n20), .A0N(\regs[12][21] ), .A1N(n20), .Y(
        n491) );
  OAI2BB2X1 U1623 ( .B0(n2212), .B1(n20), .A0N(\regs[12][22] ), .A1N(n20), .Y(
        n492) );
  OAI2BB2X1 U1624 ( .B0(n2211), .B1(n20), .A0N(\regs[12][23] ), .A1N(n20), .Y(
        n493) );
  OAI2BB2X1 U1625 ( .B0(n2210), .B1(n20), .A0N(\regs[12][24] ), .A1N(n20), .Y(
        n494) );
  OAI2BB2X1 U1626 ( .B0(n2209), .B1(n20), .A0N(\regs[12][25] ), .A1N(n20), .Y(
        n495) );
  OAI2BB2X1 U1627 ( .B0(n2208), .B1(n20), .A0N(\regs[12][26] ), .A1N(n20), .Y(
        n496) );
  OAI2BB2X1 U1628 ( .B0(n2207), .B1(n20), .A0N(\regs[12][27] ), .A1N(n20), .Y(
        n497) );
  OAI2BB2X1 U1629 ( .B0(n2206), .B1(n20), .A0N(\regs[12][28] ), .A1N(n20), .Y(
        n498) );
  OAI2BB2X1 U1630 ( .B0(n2205), .B1(n20), .A0N(\regs[12][29] ), .A1N(n20), .Y(
        n499) );
  OAI2BB2X1 U1631 ( .B0(n2204), .B1(n20), .A0N(\regs[12][30] ), .A1N(n20), .Y(
        n500) );
  OAI2BB2X1 U1632 ( .B0(n34), .B1(n20), .A0N(\regs[12][31] ), .A1N(n20), .Y(
        n501) );
  OAI2BB2X1 U1633 ( .B0(n2227), .B1(n21), .A0N(\regs[13][0] ), .A1N(n21), .Y(
        n502) );
  OAI2BB2X1 U1634 ( .B0(n2226), .B1(n21), .A0N(\regs[13][1] ), .A1N(n21), .Y(
        n503) );
  OAI2BB2X1 U1635 ( .B0(n2225), .B1(n21), .A0N(\regs[13][2] ), .A1N(n21), .Y(
        n504) );
  OAI2BB2X1 U1636 ( .B0(n6), .B1(n21), .A0N(\regs[13][3] ), .A1N(n21), .Y(n505) );
  OAI2BB2X1 U1637 ( .B0(n7), .B1(n21), .A0N(\regs[13][4] ), .A1N(n21), .Y(n506) );
  OAI2BB2X1 U1638 ( .B0(n8), .B1(n21), .A0N(\regs[13][5] ), .A1N(n21), .Y(n507) );
  OAI2BB2X1 U1639 ( .B0(n9), .B1(n21), .A0N(\regs[13][6] ), .A1N(n21), .Y(n508) );
  OAI2BB2X1 U1640 ( .B0(n2221), .B1(n21), .A0N(\regs[13][13] ), .A1N(n21), .Y(
        n515) );
  OAI2BB2X1 U1641 ( .B0(n2218), .B1(n21), .A0N(\regs[13][16] ), .A1N(n21), .Y(
        n518) );
  OAI2BB2X1 U1642 ( .B0(n2217), .B1(n21), .A0N(\regs[13][17] ), .A1N(n21), .Y(
        n519) );
  OAI2BB2X1 U1643 ( .B0(n2216), .B1(n21), .A0N(\regs[13][18] ), .A1N(n21), .Y(
        n520) );
  OAI2BB2X1 U1644 ( .B0(n2215), .B1(n21), .A0N(\regs[13][19] ), .A1N(n21), .Y(
        n521) );
  OAI2BB2X1 U1645 ( .B0(n2214), .B1(n21), .A0N(\regs[13][20] ), .A1N(n21), .Y(
        n522) );
  OAI2BB2X1 U1646 ( .B0(n2213), .B1(n21), .A0N(\regs[13][21] ), .A1N(n21), .Y(
        n523) );
  OAI2BB2X1 U1647 ( .B0(n2212), .B1(n21), .A0N(\regs[13][22] ), .A1N(n21), .Y(
        n524) );
  OAI2BB2X1 U1648 ( .B0(n2211), .B1(n21), .A0N(\regs[13][23] ), .A1N(n21), .Y(
        n525) );
  OAI2BB2X1 U1649 ( .B0(n2210), .B1(n21), .A0N(\regs[13][24] ), .A1N(n21), .Y(
        n526) );
  OAI2BB2X1 U1650 ( .B0(n2209), .B1(n21), .A0N(\regs[13][25] ), .A1N(n21), .Y(
        n527) );
  OAI2BB2X1 U1651 ( .B0(n2208), .B1(n21), .A0N(\regs[13][26] ), .A1N(n21), .Y(
        n528) );
  OAI2BB2X1 U1652 ( .B0(n2207), .B1(n21), .A0N(\regs[13][27] ), .A1N(n21), .Y(
        n529) );
  OAI2BB2X1 U1653 ( .B0(n2206), .B1(n21), .A0N(\regs[13][28] ), .A1N(n21), .Y(
        n530) );
  OAI2BB2X1 U1654 ( .B0(n2205), .B1(n21), .A0N(\regs[13][29] ), .A1N(n21), .Y(
        n531) );
  OAI2BB2X1 U1655 ( .B0(n2204), .B1(n21), .A0N(\regs[13][30] ), .A1N(n21), .Y(
        n532) );
  OAI2BB2X1 U1656 ( .B0(n34), .B1(n21), .A0N(\regs[13][31] ), .A1N(n21), .Y(
        n533) );
  OAI2BB2X1 U1657 ( .B0(n2227), .B1(n24), .A0N(\regs[14][0] ), .A1N(n24), .Y(
        n534) );
  OAI2BB2X1 U1658 ( .B0(n2226), .B1(n24), .A0N(\regs[14][1] ), .A1N(n24), .Y(
        n535) );
  OAI2BB2X1 U1659 ( .B0(n2225), .B1(n24), .A0N(\regs[14][2] ), .A1N(n24), .Y(
        n536) );
  OAI2BB2X1 U1660 ( .B0(n6), .B1(n24), .A0N(\regs[14][3] ), .A1N(n24), .Y(n537) );
  OAI2BB2X1 U1661 ( .B0(n7), .B1(n24), .A0N(\regs[14][4] ), .A1N(n24), .Y(n538) );
  OAI2BB2X1 U1662 ( .B0(n8), .B1(n24), .A0N(\regs[14][5] ), .A1N(n24), .Y(n539) );
  OAI2BB2X1 U1663 ( .B0(n9), .B1(n24), .A0N(\regs[14][6] ), .A1N(n24), .Y(n540) );
  OAI2BB2X1 U1664 ( .B0(n2221), .B1(n24), .A0N(\regs[14][13] ), .A1N(n24), .Y(
        n547) );
  OAI2BB2X1 U1665 ( .B0(n2218), .B1(n24), .A0N(\regs[14][16] ), .A1N(n24), .Y(
        n550) );
  OAI2BB2X1 U1666 ( .B0(n2217), .B1(n24), .A0N(\regs[14][17] ), .A1N(n24), .Y(
        n551) );
  OAI2BB2X1 U1667 ( .B0(n2216), .B1(n24), .A0N(\regs[14][18] ), .A1N(n24), .Y(
        n552) );
  OAI2BB2X1 U1668 ( .B0(n2215), .B1(n24), .A0N(\regs[14][19] ), .A1N(n24), .Y(
        n553) );
  OAI2BB2X1 U1669 ( .B0(n2214), .B1(n24), .A0N(\regs[14][20] ), .A1N(n24), .Y(
        n554) );
  OAI2BB2X1 U1670 ( .B0(n2213), .B1(n24), .A0N(\regs[14][21] ), .A1N(n24), .Y(
        n555) );
  OAI2BB2X1 U1671 ( .B0(n2212), .B1(n24), .A0N(\regs[14][22] ), .A1N(n24), .Y(
        n556) );
  OAI2BB2X1 U1672 ( .B0(n2211), .B1(n24), .A0N(\regs[14][23] ), .A1N(n24), .Y(
        n557) );
  OAI2BB2X1 U1673 ( .B0(n2210), .B1(n24), .A0N(\regs[14][24] ), .A1N(n24), .Y(
        n558) );
  OAI2BB2X1 U1674 ( .B0(n2209), .B1(n24), .A0N(\regs[14][25] ), .A1N(n24), .Y(
        n559) );
  OAI2BB2X1 U1675 ( .B0(n2208), .B1(n24), .A0N(\regs[14][26] ), .A1N(n24), .Y(
        n560) );
  OAI2BB2X1 U1676 ( .B0(n2207), .B1(n24), .A0N(\regs[14][27] ), .A1N(n24), .Y(
        n561) );
  OAI2BB2X1 U1677 ( .B0(n2206), .B1(n24), .A0N(\regs[14][28] ), .A1N(n24), .Y(
        n562) );
  OAI2BB2X1 U1678 ( .B0(n2205), .B1(n24), .A0N(\regs[14][29] ), .A1N(n24), .Y(
        n563) );
  OAI2BB2X1 U1679 ( .B0(n2204), .B1(n24), .A0N(\regs[14][30] ), .A1N(n24), .Y(
        n564) );
  OAI2BB2X1 U1680 ( .B0(n34), .B1(n24), .A0N(\regs[14][31] ), .A1N(n24), .Y(
        n565) );
  OAI2BB2X1 U1681 ( .B0(n2227), .B1(n61), .A0N(\regs[15][0] ), .A1N(n61), .Y(
        n566) );
  OAI2BB2X1 U1682 ( .B0(n2226), .B1(n61), .A0N(\regs[15][1] ), .A1N(n61), .Y(
        n567) );
  OAI2BB2X1 U1683 ( .B0(n2225), .B1(n61), .A0N(\regs[15][2] ), .A1N(n61), .Y(
        n568) );
  OAI2BB2X1 U1684 ( .B0(n6), .B1(n61), .A0N(\regs[15][3] ), .A1N(n61), .Y(n569) );
  OAI2BB2X1 U1685 ( .B0(n7), .B1(n61), .A0N(\regs[15][4] ), .A1N(n61), .Y(n570) );
  OAI2BB2X1 U1686 ( .B0(n8), .B1(n61), .A0N(\regs[15][5] ), .A1N(n61), .Y(n571) );
  OAI2BB2X1 U1687 ( .B0(n9), .B1(n61), .A0N(\regs[15][6] ), .A1N(n61), .Y(n572) );
  OAI2BB2X1 U1688 ( .B0(n2221), .B1(n61), .A0N(\regs[15][13] ), .A1N(n61), .Y(
        n579) );
  OAI2BB2X1 U1689 ( .B0(n2218), .B1(n61), .A0N(\regs[15][16] ), .A1N(n61), .Y(
        n582) );
  OAI2BB2X1 U1690 ( .B0(n2217), .B1(n61), .A0N(\regs[15][17] ), .A1N(n61), .Y(
        n583) );
  OAI2BB2X1 U1691 ( .B0(n2216), .B1(n61), .A0N(\regs[15][18] ), .A1N(n61), .Y(
        n584) );
  OAI2BB2X1 U1692 ( .B0(n2215), .B1(n61), .A0N(\regs[15][19] ), .A1N(n61), .Y(
        n585) );
  OAI2BB2X1 U1693 ( .B0(n2214), .B1(n61), .A0N(\regs[15][20] ), .A1N(n61), .Y(
        n586) );
  OAI2BB2X1 U1694 ( .B0(n2213), .B1(n61), .A0N(\regs[15][21] ), .A1N(n61), .Y(
        n587) );
  OAI2BB2X1 U1695 ( .B0(n2212), .B1(n61), .A0N(\regs[15][22] ), .A1N(n61), .Y(
        n588) );
  OAI2BB2X1 U1696 ( .B0(n2211), .B1(n61), .A0N(\regs[15][23] ), .A1N(n61), .Y(
        n589) );
  OAI2BB2X1 U1697 ( .B0(n2210), .B1(n61), .A0N(\regs[15][24] ), .A1N(n61), .Y(
        n590) );
  OAI2BB2X1 U1698 ( .B0(n2209), .B1(n61), .A0N(\regs[15][25] ), .A1N(n61), .Y(
        n591) );
  OAI2BB2X1 U1699 ( .B0(n2208), .B1(n61), .A0N(\regs[15][26] ), .A1N(n61), .Y(
        n592) );
  OAI2BB2X1 U1700 ( .B0(n2207), .B1(n61), .A0N(\regs[15][27] ), .A1N(n61), .Y(
        n593) );
  OAI2BB2X1 U1701 ( .B0(n2206), .B1(n61), .A0N(\regs[15][28] ), .A1N(n61), .Y(
        n594) );
  OAI2BB2X1 U1702 ( .B0(n2205), .B1(n61), .A0N(\regs[15][29] ), .A1N(n61), .Y(
        n595) );
  OAI2BB2X1 U1703 ( .B0(n2204), .B1(n61), .A0N(\regs[15][30] ), .A1N(n61), .Y(
        n596) );
  OAI2BB2X1 U1704 ( .B0(n34), .B1(n61), .A0N(\regs[15][31] ), .A1N(n61), .Y(
        n597) );
  OAI2BB2X1 U1705 ( .B0(n2227), .B1(n22), .A0N(\regs[16][0] ), .A1N(n22), .Y(
        n598) );
  OAI2BB2X1 U1706 ( .B0(n2226), .B1(n22), .A0N(\regs[16][1] ), .A1N(n22), .Y(
        n599) );
  OAI2BB2X1 U1707 ( .B0(n2225), .B1(n22), .A0N(\regs[16][2] ), .A1N(n22), .Y(
        n600) );
  OAI2BB2X1 U1708 ( .B0(n6), .B1(n22), .A0N(\regs[16][3] ), .A1N(n22), .Y(n601) );
  OAI2BB2X1 U1709 ( .B0(n7), .B1(n22), .A0N(\regs[16][4] ), .A1N(n22), .Y(n602) );
  OAI2BB2X1 U1710 ( .B0(n8), .B1(n22), .A0N(\regs[16][5] ), .A1N(n22), .Y(n603) );
  OAI2BB2X1 U1711 ( .B0(n9), .B1(n22), .A0N(\regs[16][6] ), .A1N(n22), .Y(n604) );
  OAI2BB2X1 U1712 ( .B0(n2221), .B1(n22), .A0N(\regs[16][13] ), .A1N(n22), .Y(
        n611) );
  OAI2BB2X1 U1713 ( .B0(n2218), .B1(n22), .A0N(\regs[16][16] ), .A1N(n22), .Y(
        n614) );
  OAI2BB2X1 U1714 ( .B0(n2217), .B1(n22), .A0N(\regs[16][17] ), .A1N(n22), .Y(
        n615) );
  OAI2BB2X1 U1715 ( .B0(n2216), .B1(n22), .A0N(\regs[16][18] ), .A1N(n22), .Y(
        n616) );
  OAI2BB2X1 U1716 ( .B0(n2215), .B1(n22), .A0N(\regs[16][19] ), .A1N(n22), .Y(
        n617) );
  OAI2BB2X1 U1717 ( .B0(n2214), .B1(n22), .A0N(\regs[16][20] ), .A1N(n22), .Y(
        n618) );
  OAI2BB2X1 U1718 ( .B0(n2213), .B1(n22), .A0N(\regs[16][21] ), .A1N(n22), .Y(
        n619) );
  OAI2BB2X1 U1719 ( .B0(n2212), .B1(n22), .A0N(\regs[16][22] ), .A1N(n22), .Y(
        n620) );
  OAI2BB2X1 U1720 ( .B0(n2211), .B1(n22), .A0N(\regs[16][23] ), .A1N(n22), .Y(
        n621) );
  OAI2BB2X1 U1721 ( .B0(n2210), .B1(n22), .A0N(\regs[16][24] ), .A1N(n22), .Y(
        n622) );
  OAI2BB2X1 U1722 ( .B0(n2209), .B1(n22), .A0N(\regs[16][25] ), .A1N(n22), .Y(
        n623) );
  OAI2BB2X1 U1723 ( .B0(n2208), .B1(n22), .A0N(\regs[16][26] ), .A1N(n22), .Y(
        n624) );
  OAI2BB2X1 U1724 ( .B0(n2207), .B1(n22), .A0N(\regs[16][27] ), .A1N(n22), .Y(
        n625) );
  OAI2BB2X1 U1725 ( .B0(n2206), .B1(n22), .A0N(\regs[16][28] ), .A1N(n22), .Y(
        n626) );
  OAI2BB2X1 U1726 ( .B0(n2205), .B1(n22), .A0N(\regs[16][29] ), .A1N(n22), .Y(
        n627) );
  OAI2BB2X1 U1727 ( .B0(n2204), .B1(n22), .A0N(\regs[16][30] ), .A1N(n22), .Y(
        n628) );
  OAI2BB2X1 U1728 ( .B0(n34), .B1(n22), .A0N(\regs[16][31] ), .A1N(n22), .Y(
        n629) );
  OAI2BB2X1 U1729 ( .B0(n2227), .B1(n23), .A0N(\regs[17][0] ), .A1N(n23), .Y(
        n630) );
  OAI2BB2X1 U1730 ( .B0(n2226), .B1(n23), .A0N(\regs[17][1] ), .A1N(n23), .Y(
        n631) );
  OAI2BB2X1 U1731 ( .B0(n2225), .B1(n23), .A0N(\regs[17][2] ), .A1N(n23), .Y(
        n632) );
  OAI2BB2X1 U1732 ( .B0(n6), .B1(n23), .A0N(\regs[17][3] ), .A1N(n23), .Y(n633) );
  OAI2BB2X1 U1733 ( .B0(n7), .B1(n23), .A0N(\regs[17][4] ), .A1N(n23), .Y(n634) );
  OAI2BB2X1 U1734 ( .B0(n8), .B1(n23), .A0N(\regs[17][5] ), .A1N(n23), .Y(n635) );
  OAI2BB2X1 U1735 ( .B0(n9), .B1(n23), .A0N(\regs[17][6] ), .A1N(n23), .Y(n636) );
  OAI2BB2X1 U1736 ( .B0(n2221), .B1(n23), .A0N(\regs[17][13] ), .A1N(n23), .Y(
        n643) );
  OAI2BB2X1 U1737 ( .B0(n2218), .B1(n23), .A0N(\regs[17][16] ), .A1N(n23), .Y(
        n646) );
  OAI2BB2X1 U1738 ( .B0(n2217), .B1(n23), .A0N(\regs[17][17] ), .A1N(n23), .Y(
        n647) );
  OAI2BB2X1 U1739 ( .B0(n2216), .B1(n23), .A0N(\regs[17][18] ), .A1N(n23), .Y(
        n648) );
  OAI2BB2X1 U1740 ( .B0(n2215), .B1(n23), .A0N(\regs[17][19] ), .A1N(n23), .Y(
        n649) );
  OAI2BB2X1 U1741 ( .B0(n2214), .B1(n23), .A0N(\regs[17][20] ), .A1N(n23), .Y(
        n650) );
  OAI2BB2X1 U1742 ( .B0(n2213), .B1(n23), .A0N(\regs[17][21] ), .A1N(n23), .Y(
        n651) );
  OAI2BB2X1 U1743 ( .B0(n2212), .B1(n23), .A0N(\regs[17][22] ), .A1N(n23), .Y(
        n652) );
  OAI2BB2X1 U1744 ( .B0(n2211), .B1(n23), .A0N(\regs[17][23] ), .A1N(n23), .Y(
        n653) );
  OAI2BB2X1 U1745 ( .B0(n2210), .B1(n23), .A0N(\regs[17][24] ), .A1N(n23), .Y(
        n654) );
  OAI2BB2X1 U1746 ( .B0(n2209), .B1(n23), .A0N(\regs[17][25] ), .A1N(n23), .Y(
        n655) );
  OAI2BB2X1 U1747 ( .B0(n2208), .B1(n23), .A0N(\regs[17][26] ), .A1N(n23), .Y(
        n656) );
  OAI2BB2X1 U1748 ( .B0(n2207), .B1(n23), .A0N(\regs[17][27] ), .A1N(n23), .Y(
        n657) );
  OAI2BB2X1 U1749 ( .B0(n2206), .B1(n23), .A0N(\regs[17][28] ), .A1N(n23), .Y(
        n658) );
  OAI2BB2X1 U1750 ( .B0(n2205), .B1(n23), .A0N(\regs[17][29] ), .A1N(n23), .Y(
        n659) );
  OAI2BB2X1 U1751 ( .B0(n2204), .B1(n23), .A0N(\regs[17][30] ), .A1N(n23), .Y(
        n660) );
  OAI2BB2X1 U1752 ( .B0(n34), .B1(n23), .A0N(\regs[17][31] ), .A1N(n23), .Y(
        n661) );
  OAI2BB2X1 U1753 ( .B0(n2227), .B1(n66), .A0N(\regs[18][0] ), .A1N(n66), .Y(
        n662) );
  OAI2BB2X1 U1754 ( .B0(n2226), .B1(n66), .A0N(\regs[18][1] ), .A1N(n66), .Y(
        n663) );
  OAI2BB2X1 U1755 ( .B0(n2225), .B1(n66), .A0N(\regs[18][2] ), .A1N(n66), .Y(
        n664) );
  OAI2BB2X1 U1756 ( .B0(n6), .B1(n66), .A0N(\regs[18][3] ), .A1N(n66), .Y(n665) );
  OAI2BB2X1 U1757 ( .B0(n7), .B1(n66), .A0N(\regs[18][4] ), .A1N(n66), .Y(n666) );
  OAI2BB2X1 U1758 ( .B0(n8), .B1(n66), .A0N(\regs[18][5] ), .A1N(n66), .Y(n667) );
  OAI2BB2X1 U1759 ( .B0(n9), .B1(n66), .A0N(\regs[18][6] ), .A1N(n66), .Y(n668) );
  OAI2BB2X1 U1760 ( .B0(n2221), .B1(n66), .A0N(\regs[18][13] ), .A1N(n66), .Y(
        n675) );
  OAI2BB2X1 U1761 ( .B0(n2218), .B1(n66), .A0N(\regs[18][16] ), .A1N(n66), .Y(
        n678) );
  OAI2BB2X1 U1762 ( .B0(n2217), .B1(n66), .A0N(\regs[18][17] ), .A1N(n66), .Y(
        n679) );
  OAI2BB2X1 U1763 ( .B0(n2216), .B1(n66), .A0N(\regs[18][18] ), .A1N(n66), .Y(
        n680) );
  OAI2BB2X1 U1764 ( .B0(n2215), .B1(n66), .A0N(\regs[18][19] ), .A1N(n66), .Y(
        n681) );
  OAI2BB2X1 U1765 ( .B0(n2214), .B1(n66), .A0N(\regs[18][20] ), .A1N(n66), .Y(
        n682) );
  OAI2BB2X1 U1766 ( .B0(n2213), .B1(n66), .A0N(\regs[18][21] ), .A1N(n66), .Y(
        n683) );
  OAI2BB2X1 U1767 ( .B0(n2212), .B1(n66), .A0N(\regs[18][22] ), .A1N(n66), .Y(
        n684) );
  OAI2BB2X1 U1768 ( .B0(n2211), .B1(n66), .A0N(\regs[18][23] ), .A1N(n66), .Y(
        n685) );
  OAI2BB2X1 U1769 ( .B0(n2210), .B1(n66), .A0N(\regs[18][24] ), .A1N(n66), .Y(
        n686) );
  OAI2BB2X1 U1770 ( .B0(n2209), .B1(n66), .A0N(\regs[18][25] ), .A1N(n66), .Y(
        n687) );
  OAI2BB2X1 U1771 ( .B0(n2208), .B1(n66), .A0N(\regs[18][26] ), .A1N(n66), .Y(
        n688) );
  OAI2BB2X1 U1772 ( .B0(n2207), .B1(n66), .A0N(\regs[18][27] ), .A1N(n66), .Y(
        n689) );
  OAI2BB2X1 U1773 ( .B0(n2206), .B1(n66), .A0N(\regs[18][28] ), .A1N(n66), .Y(
        n690) );
  OAI2BB2X1 U1774 ( .B0(n2205), .B1(n66), .A0N(\regs[18][29] ), .A1N(n66), .Y(
        n691) );
  OAI2BB2X1 U1775 ( .B0(n2204), .B1(n66), .A0N(\regs[18][30] ), .A1N(n66), .Y(
        n692) );
  OAI2BB2X1 U1776 ( .B0(n34), .B1(n66), .A0N(\regs[18][31] ), .A1N(n66), .Y(
        n693) );
  OAI2BB2X1 U1777 ( .B0(n2227), .B1(n67), .A0N(\regs[19][0] ), .A1N(n67), .Y(
        n694) );
  OAI2BB2X1 U1778 ( .B0(n2226), .B1(n67), .A0N(\regs[19][1] ), .A1N(n67), .Y(
        n695) );
  OAI2BB2X1 U1779 ( .B0(n2225), .B1(n67), .A0N(\regs[19][2] ), .A1N(n67), .Y(
        n696) );
  OAI2BB2X1 U1780 ( .B0(n6), .B1(n67), .A0N(\regs[19][3] ), .A1N(n67), .Y(n697) );
  OAI2BB2X1 U1781 ( .B0(n7), .B1(n67), .A0N(\regs[19][4] ), .A1N(n67), .Y(n698) );
  OAI2BB2X1 U1782 ( .B0(n8), .B1(n67), .A0N(\regs[19][5] ), .A1N(n67), .Y(n699) );
  OAI2BB2X1 U1783 ( .B0(n9), .B1(n67), .A0N(\regs[19][6] ), .A1N(n67), .Y(n700) );
  OAI2BB2X1 U1784 ( .B0(n2221), .B1(n67), .A0N(\regs[19][13] ), .A1N(n67), .Y(
        n707) );
  OAI2BB2X1 U1785 ( .B0(n2218), .B1(n67), .A0N(\regs[19][16] ), .A1N(n67), .Y(
        n710) );
  OAI2BB2X1 U1786 ( .B0(n2217), .B1(n67), .A0N(\regs[19][17] ), .A1N(n67), .Y(
        n711) );
  OAI2BB2X1 U1787 ( .B0(n2216), .B1(n67), .A0N(\regs[19][18] ), .A1N(n67), .Y(
        n712) );
  OAI2BB2X1 U1788 ( .B0(n2215), .B1(n67), .A0N(\regs[19][19] ), .A1N(n67), .Y(
        n713) );
  OAI2BB2X1 U1789 ( .B0(n2214), .B1(n67), .A0N(\regs[19][20] ), .A1N(n67), .Y(
        n714) );
  OAI2BB2X1 U1790 ( .B0(n2213), .B1(n67), .A0N(\regs[19][21] ), .A1N(n67), .Y(
        n715) );
  OAI2BB2X1 U1791 ( .B0(n2212), .B1(n67), .A0N(\regs[19][22] ), .A1N(n67), .Y(
        n716) );
  OAI2BB2X1 U1792 ( .B0(n2211), .B1(n67), .A0N(\regs[19][23] ), .A1N(n67), .Y(
        n717) );
  OAI2BB2X1 U1793 ( .B0(n2210), .B1(n67), .A0N(\regs[19][24] ), .A1N(n67), .Y(
        n718) );
  OAI2BB2X1 U1794 ( .B0(n2209), .B1(n67), .A0N(\regs[19][25] ), .A1N(n67), .Y(
        n719) );
  OAI2BB2X1 U1795 ( .B0(n2208), .B1(n67), .A0N(\regs[19][26] ), .A1N(n67), .Y(
        n720) );
  OAI2BB2X1 U1796 ( .B0(n2207), .B1(n67), .A0N(\regs[19][27] ), .A1N(n67), .Y(
        n721) );
  OAI2BB2X1 U1797 ( .B0(n2206), .B1(n67), .A0N(\regs[19][28] ), .A1N(n67), .Y(
        n722) );
  OAI2BB2X1 U1798 ( .B0(n2205), .B1(n67), .A0N(\regs[19][29] ), .A1N(n67), .Y(
        n723) );
  OAI2BB2X1 U1799 ( .B0(n2204), .B1(n67), .A0N(\regs[19][30] ), .A1N(n67), .Y(
        n724) );
  OAI2BB2X1 U1800 ( .B0(n34), .B1(n67), .A0N(\regs[19][31] ), .A1N(n67), .Y(
        n725) );
  OAI2BB2X1 U1801 ( .B0(n2227), .B1(n25), .A0N(\regs[20][0] ), .A1N(n25), .Y(
        n726) );
  OAI2BB2X1 U1802 ( .B0(n2226), .B1(n25), .A0N(\regs[20][1] ), .A1N(n25), .Y(
        n727) );
  OAI2BB2X1 U1803 ( .B0(n2225), .B1(n25), .A0N(\regs[20][2] ), .A1N(n25), .Y(
        n728) );
  OAI2BB2X1 U1804 ( .B0(n6), .B1(n25), .A0N(\regs[20][3] ), .A1N(n25), .Y(n729) );
  OAI2BB2X1 U1805 ( .B0(n7), .B1(n25), .A0N(\regs[20][4] ), .A1N(n25), .Y(n730) );
  OAI2BB2X1 U1806 ( .B0(n8), .B1(n25), .A0N(\regs[20][5] ), .A1N(n25), .Y(n731) );
  OAI2BB2X1 U1807 ( .B0(n9), .B1(n25), .A0N(\regs[20][6] ), .A1N(n25), .Y(n732) );
  OAI2BB2X1 U1808 ( .B0(n2221), .B1(n25), .A0N(\regs[20][13] ), .A1N(n25), .Y(
        n739) );
  OAI2BB2X1 U1809 ( .B0(n2218), .B1(n25), .A0N(\regs[20][16] ), .A1N(n25), .Y(
        n742) );
  OAI2BB2X1 U1810 ( .B0(n2217), .B1(n25), .A0N(\regs[20][17] ), .A1N(n25), .Y(
        n743) );
  OAI2BB2X1 U1811 ( .B0(n2216), .B1(n25), .A0N(\regs[20][18] ), .A1N(n25), .Y(
        n744) );
  OAI2BB2X1 U1812 ( .B0(n2215), .B1(n25), .A0N(\regs[20][19] ), .A1N(n25), .Y(
        n745) );
  OAI2BB2X1 U1813 ( .B0(n2214), .B1(n25), .A0N(\regs[20][20] ), .A1N(n25), .Y(
        n746) );
  OAI2BB2X1 U1814 ( .B0(n2213), .B1(n25), .A0N(\regs[20][21] ), .A1N(n25), .Y(
        n747) );
  OAI2BB2X1 U1815 ( .B0(n2212), .B1(n25), .A0N(\regs[20][22] ), .A1N(n25), .Y(
        n748) );
  OAI2BB2X1 U1816 ( .B0(n2211), .B1(n25), .A0N(\regs[20][23] ), .A1N(n25), .Y(
        n749) );
  OAI2BB2X1 U1817 ( .B0(n2210), .B1(n25), .A0N(\regs[20][24] ), .A1N(n25), .Y(
        n750) );
  OAI2BB2X1 U1818 ( .B0(n2209), .B1(n25), .A0N(\regs[20][25] ), .A1N(n25), .Y(
        n751) );
  OAI2BB2X1 U1819 ( .B0(n2208), .B1(n25), .A0N(\regs[20][26] ), .A1N(n25), .Y(
        n752) );
  OAI2BB2X1 U1820 ( .B0(n2207), .B1(n25), .A0N(\regs[20][27] ), .A1N(n25), .Y(
        n753) );
  OAI2BB2X1 U1821 ( .B0(n2206), .B1(n25), .A0N(\regs[20][28] ), .A1N(n25), .Y(
        n754) );
  OAI2BB2X1 U1822 ( .B0(n2205), .B1(n25), .A0N(\regs[20][29] ), .A1N(n25), .Y(
        n755) );
  OAI2BB2X1 U1823 ( .B0(n2204), .B1(n25), .A0N(\regs[20][30] ), .A1N(n25), .Y(
        n756) );
  OAI2BB2X1 U1824 ( .B0(n34), .B1(n25), .A0N(\regs[20][31] ), .A1N(n25), .Y(
        n757) );
  OAI2BB2X1 U1825 ( .B0(n2227), .B1(n26), .A0N(\regs[21][0] ), .A1N(n26), .Y(
        n758) );
  OAI2BB2X1 U1826 ( .B0(n2226), .B1(n26), .A0N(\regs[21][1] ), .A1N(n26), .Y(
        n759) );
  OAI2BB2X1 U1827 ( .B0(n2225), .B1(n26), .A0N(\regs[21][2] ), .A1N(n26), .Y(
        n760) );
  OAI2BB2X1 U1828 ( .B0(n6), .B1(n26), .A0N(\regs[21][3] ), .A1N(n26), .Y(n761) );
  OAI2BB2X1 U1829 ( .B0(n7), .B1(n26), .A0N(\regs[21][4] ), .A1N(n26), .Y(n762) );
  OAI2BB2X1 U1830 ( .B0(n8), .B1(n26), .A0N(\regs[21][5] ), .A1N(n26), .Y(n763) );
  OAI2BB2X1 U1831 ( .B0(n9), .B1(n26), .A0N(\regs[21][6] ), .A1N(n26), .Y(n764) );
  OAI2BB2X1 U1832 ( .B0(n2221), .B1(n26), .A0N(\regs[21][13] ), .A1N(n26), .Y(
        n771) );
  OAI2BB2X1 U1833 ( .B0(n2218), .B1(n26), .A0N(\regs[21][16] ), .A1N(n26), .Y(
        n774) );
  OAI2BB2X1 U1834 ( .B0(n2217), .B1(n26), .A0N(\regs[21][17] ), .A1N(n26), .Y(
        n775) );
  OAI2BB2X1 U1835 ( .B0(n2216), .B1(n26), .A0N(\regs[21][18] ), .A1N(n26), .Y(
        n776) );
  OAI2BB2X1 U1836 ( .B0(n2215), .B1(n26), .A0N(\regs[21][19] ), .A1N(n26), .Y(
        n777) );
  OAI2BB2X1 U1837 ( .B0(n2214), .B1(n26), .A0N(\regs[21][20] ), .A1N(n26), .Y(
        n778) );
  OAI2BB2X1 U1838 ( .B0(n2213), .B1(n26), .A0N(\regs[21][21] ), .A1N(n26), .Y(
        n779) );
  OAI2BB2X1 U1839 ( .B0(n2212), .B1(n26), .A0N(\regs[21][22] ), .A1N(n26), .Y(
        n780) );
  OAI2BB2X1 U1840 ( .B0(n2211), .B1(n26), .A0N(\regs[21][23] ), .A1N(n26), .Y(
        n781) );
  OAI2BB2X1 U1841 ( .B0(n2210), .B1(n26), .A0N(\regs[21][24] ), .A1N(n26), .Y(
        n782) );
  OAI2BB2X1 U1842 ( .B0(n2209), .B1(n26), .A0N(\regs[21][25] ), .A1N(n26), .Y(
        n783) );
  OAI2BB2X1 U1843 ( .B0(n2208), .B1(n26), .A0N(\regs[21][26] ), .A1N(n26), .Y(
        n784) );
  OAI2BB2X1 U1844 ( .B0(n2207), .B1(n26), .A0N(\regs[21][27] ), .A1N(n26), .Y(
        n785) );
  OAI2BB2X1 U1845 ( .B0(n2206), .B1(n26), .A0N(\regs[21][28] ), .A1N(n26), .Y(
        n786) );
  OAI2BB2X1 U1846 ( .B0(n2205), .B1(n26), .A0N(\regs[21][29] ), .A1N(n26), .Y(
        n787) );
  OAI2BB2X1 U1847 ( .B0(n2204), .B1(n26), .A0N(\regs[21][30] ), .A1N(n26), .Y(
        n788) );
  OAI2BB2X1 U1848 ( .B0(n34), .B1(n26), .A0N(\regs[21][31] ), .A1N(n26), .Y(
        n789) );
  OAI2BB2X1 U1849 ( .B0(n2227), .B1(n27), .A0N(\regs[22][0] ), .A1N(n27), .Y(
        n790) );
  OAI2BB2X1 U1850 ( .B0(n2226), .B1(n27), .A0N(\regs[22][1] ), .A1N(n27), .Y(
        n791) );
  OAI2BB2X1 U1851 ( .B0(n2225), .B1(n27), .A0N(\regs[22][2] ), .A1N(n27), .Y(
        n792) );
  OAI2BB2X1 U1852 ( .B0(n6), .B1(n27), .A0N(\regs[22][3] ), .A1N(n27), .Y(n793) );
  OAI2BB2X1 U1853 ( .B0(n7), .B1(n27), .A0N(\regs[22][4] ), .A1N(n27), .Y(n794) );
  OAI2BB2X1 U1854 ( .B0(n8), .B1(n27), .A0N(\regs[22][5] ), .A1N(n27), .Y(n795) );
  OAI2BB2X1 U1855 ( .B0(n9), .B1(n27), .A0N(\regs[22][6] ), .A1N(n27), .Y(n796) );
  OAI2BB2X1 U1856 ( .B0(n2221), .B1(n27), .A0N(\regs[22][13] ), .A1N(n27), .Y(
        n803) );
  OAI2BB2X1 U1857 ( .B0(n2218), .B1(n27), .A0N(\regs[22][16] ), .A1N(n27), .Y(
        n806) );
  OAI2BB2X1 U1858 ( .B0(n2217), .B1(n27), .A0N(\regs[22][17] ), .A1N(n27), .Y(
        n807) );
  OAI2BB2X1 U1859 ( .B0(n2216), .B1(n27), .A0N(\regs[22][18] ), .A1N(n27), .Y(
        n808) );
  OAI2BB2X1 U1860 ( .B0(n2215), .B1(n27), .A0N(\regs[22][19] ), .A1N(n27), .Y(
        n809) );
  OAI2BB2X1 U1861 ( .B0(n2214), .B1(n27), .A0N(\regs[22][20] ), .A1N(n27), .Y(
        n810) );
  OAI2BB2X1 U1862 ( .B0(n2213), .B1(n27), .A0N(\regs[22][21] ), .A1N(n27), .Y(
        n811) );
  OAI2BB2X1 U1863 ( .B0(n2212), .B1(n27), .A0N(\regs[22][22] ), .A1N(n27), .Y(
        n812) );
  OAI2BB2X1 U1864 ( .B0(n2211), .B1(n27), .A0N(\regs[22][23] ), .A1N(n27), .Y(
        n813) );
  OAI2BB2X1 U1865 ( .B0(n2210), .B1(n27), .A0N(\regs[22][24] ), .A1N(n27), .Y(
        n814) );
  OAI2BB2X1 U1866 ( .B0(n2209), .B1(n27), .A0N(\regs[22][25] ), .A1N(n27), .Y(
        n815) );
  OAI2BB2X1 U1867 ( .B0(n2208), .B1(n27), .A0N(\regs[22][26] ), .A1N(n27), .Y(
        n816) );
  OAI2BB2X1 U1868 ( .B0(n2207), .B1(n27), .A0N(\regs[22][27] ), .A1N(n27), .Y(
        n817) );
  OAI2BB2X1 U1869 ( .B0(n2206), .B1(n27), .A0N(\regs[22][28] ), .A1N(n27), .Y(
        n818) );
  OAI2BB2X1 U1870 ( .B0(n2205), .B1(n27), .A0N(\regs[22][29] ), .A1N(n27), .Y(
        n819) );
  OAI2BB2X1 U1871 ( .B0(n2204), .B1(n27), .A0N(\regs[22][30] ), .A1N(n27), .Y(
        n820) );
  OAI2BB2X1 U1872 ( .B0(n34), .B1(n27), .A0N(\regs[22][31] ), .A1N(n27), .Y(
        n821) );
  OAI2BB2X1 U1873 ( .B0(n2227), .B1(n28), .A0N(\regs[23][0] ), .A1N(n28), .Y(
        n822) );
  OAI2BB2X1 U1874 ( .B0(n2226), .B1(n28), .A0N(\regs[23][1] ), .A1N(n28), .Y(
        n823) );
  OAI2BB2X1 U1875 ( .B0(n2225), .B1(n28), .A0N(\regs[23][2] ), .A1N(n28), .Y(
        n824) );
  OAI2BB2X1 U1876 ( .B0(n6), .B1(n28), .A0N(\regs[23][3] ), .A1N(n28), .Y(n825) );
  OAI2BB2X1 U1877 ( .B0(n7), .B1(n28), .A0N(\regs[23][4] ), .A1N(n28), .Y(n826) );
  OAI2BB2X1 U1878 ( .B0(n8), .B1(n28), .A0N(\regs[23][5] ), .A1N(n28), .Y(n827) );
  OAI2BB2X1 U1879 ( .B0(n9), .B1(n28), .A0N(\regs[23][6] ), .A1N(n28), .Y(n828) );
  OAI2BB2X1 U1880 ( .B0(n2221), .B1(n28), .A0N(\regs[23][13] ), .A1N(n28), .Y(
        n835) );
  OAI2BB2X1 U1881 ( .B0(n2218), .B1(n28), .A0N(\regs[23][16] ), .A1N(n28), .Y(
        n838) );
  OAI2BB2X1 U1882 ( .B0(n2217), .B1(n28), .A0N(\regs[23][17] ), .A1N(n28), .Y(
        n839) );
  OAI2BB2X1 U1883 ( .B0(n2216), .B1(n28), .A0N(\regs[23][18] ), .A1N(n28), .Y(
        n840) );
  OAI2BB2X1 U1884 ( .B0(n2215), .B1(n28), .A0N(\regs[23][19] ), .A1N(n28), .Y(
        n841) );
  OAI2BB2X1 U1885 ( .B0(n2214), .B1(n28), .A0N(\regs[23][20] ), .A1N(n28), .Y(
        n842) );
  OAI2BB2X1 U1886 ( .B0(n2213), .B1(n28), .A0N(\regs[23][21] ), .A1N(n28), .Y(
        n843) );
  OAI2BB2X1 U1887 ( .B0(n2212), .B1(n28), .A0N(\regs[23][22] ), .A1N(n28), .Y(
        n844) );
  OAI2BB2X1 U1888 ( .B0(n2211), .B1(n28), .A0N(\regs[23][23] ), .A1N(n28), .Y(
        n845) );
  OAI2BB2X1 U1889 ( .B0(n2210), .B1(n28), .A0N(\regs[23][24] ), .A1N(n28), .Y(
        n846) );
  OAI2BB2X1 U1890 ( .B0(n2209), .B1(n28), .A0N(\regs[23][25] ), .A1N(n28), .Y(
        n847) );
  OAI2BB2X1 U1891 ( .B0(n2208), .B1(n28), .A0N(\regs[23][26] ), .A1N(n28), .Y(
        n848) );
  OAI2BB2X1 U1892 ( .B0(n2207), .B1(n28), .A0N(\regs[23][27] ), .A1N(n28), .Y(
        n849) );
  OAI2BB2X1 U1893 ( .B0(n2206), .B1(n28), .A0N(\regs[23][28] ), .A1N(n28), .Y(
        n850) );
  OAI2BB2X1 U1894 ( .B0(n2205), .B1(n28), .A0N(\regs[23][29] ), .A1N(n28), .Y(
        n851) );
  OAI2BB2X1 U1895 ( .B0(n2204), .B1(n28), .A0N(\regs[23][30] ), .A1N(n28), .Y(
        n852) );
  OAI2BB2X1 U1896 ( .B0(n34), .B1(n28), .A0N(\regs[23][31] ), .A1N(n28), .Y(
        n853) );
  OAI2BB2X1 U1897 ( .B0(n2227), .B1(n29), .A0N(\regs[24][0] ), .A1N(n29), .Y(
        n854) );
  OAI2BB2X1 U1898 ( .B0(n2226), .B1(n29), .A0N(\regs[24][1] ), .A1N(n29), .Y(
        n855) );
  OAI2BB2X1 U1899 ( .B0(n2225), .B1(n29), .A0N(\regs[24][2] ), .A1N(n29), .Y(
        n856) );
  OAI2BB2X1 U1900 ( .B0(n6), .B1(n29), .A0N(\regs[24][3] ), .A1N(n29), .Y(n857) );
  OAI2BB2X1 U1901 ( .B0(n7), .B1(n29), .A0N(\regs[24][4] ), .A1N(n29), .Y(n858) );
  OAI2BB2X1 U1902 ( .B0(n8), .B1(n29), .A0N(\regs[24][5] ), .A1N(n29), .Y(n859) );
  OAI2BB2X1 U1903 ( .B0(n9), .B1(n29), .A0N(\regs[24][6] ), .A1N(n29), .Y(n860) );
  OAI2BB2X1 U1904 ( .B0(n2221), .B1(n29), .A0N(\regs[24][13] ), .A1N(n29), .Y(
        n867) );
  OAI2BB2X1 U1905 ( .B0(n2218), .B1(n29), .A0N(\regs[24][16] ), .A1N(n29), .Y(
        n870) );
  OAI2BB2X1 U1906 ( .B0(n2217), .B1(n29), .A0N(\regs[24][17] ), .A1N(n29), .Y(
        n871) );
  OAI2BB2X1 U1907 ( .B0(n2216), .B1(n29), .A0N(\regs[24][18] ), .A1N(n29), .Y(
        n872) );
  OAI2BB2X1 U1908 ( .B0(n2215), .B1(n29), .A0N(\regs[24][19] ), .A1N(n29), .Y(
        n873) );
  OAI2BB2X1 U1909 ( .B0(n2214), .B1(n29), .A0N(\regs[24][20] ), .A1N(n29), .Y(
        n874) );
  OAI2BB2X1 U1910 ( .B0(n2213), .B1(n29), .A0N(\regs[24][21] ), .A1N(n29), .Y(
        n875) );
  OAI2BB2X1 U1911 ( .B0(n2212), .B1(n29), .A0N(\regs[24][22] ), .A1N(n29), .Y(
        n876) );
  OAI2BB2X1 U1912 ( .B0(n2211), .B1(n29), .A0N(\regs[24][23] ), .A1N(n29), .Y(
        n877) );
  OAI2BB2X1 U1913 ( .B0(n2210), .B1(n29), .A0N(\regs[24][24] ), .A1N(n29), .Y(
        n878) );
  OAI2BB2X1 U1914 ( .B0(n2209), .B1(n29), .A0N(\regs[24][25] ), .A1N(n29), .Y(
        n879) );
  OAI2BB2X1 U1915 ( .B0(n2208), .B1(n29), .A0N(\regs[24][26] ), .A1N(n29), .Y(
        n880) );
  OAI2BB2X1 U1916 ( .B0(n2207), .B1(n29), .A0N(\regs[24][27] ), .A1N(n29), .Y(
        n881) );
  OAI2BB2X1 U1917 ( .B0(n2206), .B1(n29), .A0N(\regs[24][28] ), .A1N(n29), .Y(
        n882) );
  OAI2BB2X1 U1918 ( .B0(n2205), .B1(n29), .A0N(\regs[24][29] ), .A1N(n29), .Y(
        n883) );
  OAI2BB2X1 U1919 ( .B0(n2204), .B1(n29), .A0N(\regs[24][30] ), .A1N(n29), .Y(
        n884) );
  OAI2BB2X1 U1920 ( .B0(n34), .B1(n29), .A0N(\regs[24][31] ), .A1N(n29), .Y(
        n885) );
  OAI2BB2X1 U1921 ( .B0(n2227), .B1(n30), .A0N(\regs[25][0] ), .A1N(n30), .Y(
        n886) );
  OAI2BB2X1 U1922 ( .B0(n2226), .B1(n30), .A0N(\regs[25][1] ), .A1N(n30), .Y(
        n887) );
  OAI2BB2X1 U1923 ( .B0(n2225), .B1(n30), .A0N(\regs[25][2] ), .A1N(n30), .Y(
        n888) );
  OAI2BB2X1 U1924 ( .B0(n6), .B1(n30), .A0N(\regs[25][3] ), .A1N(n30), .Y(n889) );
  OAI2BB2X1 U1925 ( .B0(n7), .B1(n30), .A0N(\regs[25][4] ), .A1N(n30), .Y(n890) );
  OAI2BB2X1 U1926 ( .B0(n8), .B1(n30), .A0N(\regs[25][5] ), .A1N(n30), .Y(n891) );
  OAI2BB2X1 U1927 ( .B0(n9), .B1(n30), .A0N(\regs[25][6] ), .A1N(n30), .Y(n892) );
  OAI2BB2X1 U1928 ( .B0(n2221), .B1(n30), .A0N(\regs[25][13] ), .A1N(n30), .Y(
        n899) );
  OAI2BB2X1 U1929 ( .B0(n2218), .B1(n30), .A0N(\regs[25][16] ), .A1N(n30), .Y(
        n902) );
  OAI2BB2X1 U1930 ( .B0(n2217), .B1(n30), .A0N(\regs[25][17] ), .A1N(n30), .Y(
        n903) );
  OAI2BB2X1 U1931 ( .B0(n2216), .B1(n30), .A0N(\regs[25][18] ), .A1N(n30), .Y(
        n904) );
  OAI2BB2X1 U1932 ( .B0(n2215), .B1(n30), .A0N(\regs[25][19] ), .A1N(n30), .Y(
        n905) );
  OAI2BB2X1 U1933 ( .B0(n2214), .B1(n30), .A0N(\regs[25][20] ), .A1N(n30), .Y(
        n906) );
  OAI2BB2X1 U1934 ( .B0(n2213), .B1(n30), .A0N(\regs[25][21] ), .A1N(n30), .Y(
        n907) );
  OAI2BB2X1 U1935 ( .B0(n2212), .B1(n30), .A0N(\regs[25][22] ), .A1N(n30), .Y(
        n908) );
  OAI2BB2X1 U1936 ( .B0(n2211), .B1(n30), .A0N(\regs[25][23] ), .A1N(n30), .Y(
        n909) );
  OAI2BB2X1 U1937 ( .B0(n2210), .B1(n30), .A0N(\regs[25][24] ), .A1N(n30), .Y(
        n910) );
  OAI2BB2X1 U1938 ( .B0(n2209), .B1(n30), .A0N(\regs[25][25] ), .A1N(n30), .Y(
        n911) );
  OAI2BB2X1 U1939 ( .B0(n2208), .B1(n30), .A0N(\regs[25][26] ), .A1N(n30), .Y(
        n912) );
  OAI2BB2X1 U1940 ( .B0(n2207), .B1(n30), .A0N(\regs[25][27] ), .A1N(n30), .Y(
        n913) );
  OAI2BB2X1 U1941 ( .B0(n2206), .B1(n30), .A0N(\regs[25][28] ), .A1N(n30), .Y(
        n914) );
  OAI2BB2X1 U1942 ( .B0(n2205), .B1(n30), .A0N(\regs[25][29] ), .A1N(n30), .Y(
        n915) );
  OAI2BB2X1 U1943 ( .B0(n2204), .B1(n30), .A0N(\regs[25][30] ), .A1N(n30), .Y(
        n916) );
  OAI2BB2X1 U1944 ( .B0(n34), .B1(n30), .A0N(\regs[25][31] ), .A1N(n30), .Y(
        n917) );
  OAI2BB2X1 U1945 ( .B0(n2227), .B1(n31), .A0N(\regs[26][0] ), .A1N(n31), .Y(
        n918) );
  OAI2BB2X1 U1946 ( .B0(n2226), .B1(n31), .A0N(\regs[26][1] ), .A1N(n31), .Y(
        n919) );
  OAI2BB2X1 U1947 ( .B0(n2225), .B1(n31), .A0N(\regs[26][2] ), .A1N(n31), .Y(
        n920) );
  OAI2BB2X1 U1948 ( .B0(n6), .B1(n31), .A0N(\regs[26][3] ), .A1N(n31), .Y(n921) );
  OAI2BB2X1 U1949 ( .B0(n7), .B1(n31), .A0N(\regs[26][4] ), .A1N(n31), .Y(n922) );
  OAI2BB2X1 U1950 ( .B0(n8), .B1(n31), .A0N(\regs[26][5] ), .A1N(n31), .Y(n923) );
  OAI2BB2X1 U1951 ( .B0(n9), .B1(n31), .A0N(\regs[26][6] ), .A1N(n31), .Y(n924) );
  OAI2BB2X1 U1952 ( .B0(n2221), .B1(n31), .A0N(\regs[26][13] ), .A1N(n31), .Y(
        n931) );
  OAI2BB2X1 U1953 ( .B0(n2218), .B1(n31), .A0N(\regs[26][16] ), .A1N(n31), .Y(
        n934) );
  OAI2BB2X1 U1954 ( .B0(n2217), .B1(n31), .A0N(\regs[26][17] ), .A1N(n31), .Y(
        n935) );
  OAI2BB2X1 U1955 ( .B0(n2216), .B1(n31), .A0N(\regs[26][18] ), .A1N(n31), .Y(
        n936) );
  OAI2BB2X1 U1956 ( .B0(n2215), .B1(n31), .A0N(\regs[26][19] ), .A1N(n31), .Y(
        n937) );
  OAI2BB2X1 U1957 ( .B0(n2214), .B1(n31), .A0N(\regs[26][20] ), .A1N(n31), .Y(
        n938) );
  OAI2BB2X1 U1958 ( .B0(n2213), .B1(n31), .A0N(\regs[26][21] ), .A1N(n31), .Y(
        n939) );
  OAI2BB2X1 U1959 ( .B0(n2212), .B1(n31), .A0N(\regs[26][22] ), .A1N(n31), .Y(
        n940) );
  OAI2BB2X1 U1960 ( .B0(n2211), .B1(n31), .A0N(\regs[26][23] ), .A1N(n31), .Y(
        n941) );
  OAI2BB2X1 U1961 ( .B0(n2210), .B1(n31), .A0N(\regs[26][24] ), .A1N(n31), .Y(
        n942) );
  OAI2BB2X1 U1962 ( .B0(n2209), .B1(n31), .A0N(\regs[26][25] ), .A1N(n31), .Y(
        n943) );
  OAI2BB2X1 U1963 ( .B0(n2208), .B1(n31), .A0N(\regs[26][26] ), .A1N(n31), .Y(
        n944) );
  OAI2BB2X1 U1964 ( .B0(n2207), .B1(n31), .A0N(\regs[26][27] ), .A1N(n31), .Y(
        n945) );
  OAI2BB2X1 U1965 ( .B0(n2206), .B1(n31), .A0N(\regs[26][28] ), .A1N(n31), .Y(
        n946) );
  OAI2BB2X1 U1966 ( .B0(n2205), .B1(n31), .A0N(\regs[26][29] ), .A1N(n31), .Y(
        n947) );
  OAI2BB2X1 U1967 ( .B0(n2204), .B1(n31), .A0N(\regs[26][30] ), .A1N(n31), .Y(
        n948) );
  OAI2BB2X1 U1968 ( .B0(n34), .B1(n31), .A0N(\regs[26][31] ), .A1N(n31), .Y(
        n949) );
  OAI2BB2X1 U1969 ( .B0(n2227), .B1(n32), .A0N(\regs[27][0] ), .A1N(n32), .Y(
        n950) );
  OAI2BB2X1 U1970 ( .B0(n2226), .B1(n32), .A0N(\regs[27][1] ), .A1N(n32), .Y(
        n951) );
  OAI2BB2X1 U1971 ( .B0(n2225), .B1(n32), .A0N(\regs[27][2] ), .A1N(n32), .Y(
        n952) );
  OAI2BB2X1 U1972 ( .B0(n6), .B1(n32), .A0N(\regs[27][3] ), .A1N(n32), .Y(n953) );
  OAI2BB2X1 U1973 ( .B0(n7), .B1(n32), .A0N(\regs[27][4] ), .A1N(n32), .Y(n954) );
  OAI2BB2X1 U1974 ( .B0(n8), .B1(n32), .A0N(\regs[27][5] ), .A1N(n32), .Y(n955) );
  OAI2BB2X1 U1975 ( .B0(n9), .B1(n32), .A0N(\regs[27][6] ), .A1N(n32), .Y(n956) );
  OAI2BB2X1 U1976 ( .B0(n2221), .B1(n32), .A0N(\regs[27][13] ), .A1N(n32), .Y(
        n963) );
  OAI2BB2X1 U1977 ( .B0(n2218), .B1(n32), .A0N(\regs[27][16] ), .A1N(n32), .Y(
        n966) );
  OAI2BB2X1 U1978 ( .B0(n2217), .B1(n32), .A0N(\regs[27][17] ), .A1N(n32), .Y(
        n967) );
  OAI2BB2X1 U1979 ( .B0(n2216), .B1(n32), .A0N(\regs[27][18] ), .A1N(n32), .Y(
        n968) );
  OAI2BB2X1 U1980 ( .B0(n2215), .B1(n32), .A0N(\regs[27][19] ), .A1N(n32), .Y(
        n969) );
  OAI2BB2X1 U1981 ( .B0(n2214), .B1(n32), .A0N(\regs[27][20] ), .A1N(n32), .Y(
        n970) );
  OAI2BB2X1 U1982 ( .B0(n2213), .B1(n32), .A0N(\regs[27][21] ), .A1N(n32), .Y(
        n971) );
  OAI2BB2X1 U1983 ( .B0(n2212), .B1(n32), .A0N(\regs[27][22] ), .A1N(n32), .Y(
        n972) );
  OAI2BB2X1 U1984 ( .B0(n2211), .B1(n32), .A0N(\regs[27][23] ), .A1N(n32), .Y(
        n973) );
  OAI2BB2X1 U1985 ( .B0(n2210), .B1(n32), .A0N(\regs[27][24] ), .A1N(n32), .Y(
        n974) );
  OAI2BB2X1 U1986 ( .B0(n2209), .B1(n32), .A0N(\regs[27][25] ), .A1N(n32), .Y(
        n975) );
  OAI2BB2X1 U1987 ( .B0(n2208), .B1(n32), .A0N(\regs[27][26] ), .A1N(n32), .Y(
        n976) );
  OAI2BB2X1 U1988 ( .B0(n2207), .B1(n32), .A0N(\regs[27][27] ), .A1N(n32), .Y(
        n977) );
  OAI2BB2X1 U1989 ( .B0(n2206), .B1(n32), .A0N(\regs[27][28] ), .A1N(n32), .Y(
        n978) );
  OAI2BB2X1 U1990 ( .B0(n2205), .B1(n32), .A0N(\regs[27][29] ), .A1N(n32), .Y(
        n979) );
  OAI2BB2X1 U1991 ( .B0(n2204), .B1(n32), .A0N(\regs[27][30] ), .A1N(n32), .Y(
        n980) );
  OAI2BB2X1 U1992 ( .B0(n34), .B1(n32), .A0N(\regs[27][31] ), .A1N(n32), .Y(
        n981) );
  OAI2BB2X1 U1993 ( .B0(n2227), .B1(n33), .A0N(\regs[28][0] ), .A1N(n33), .Y(
        n982) );
  OAI2BB2X1 U1994 ( .B0(n2226), .B1(n33), .A0N(\regs[28][1] ), .A1N(n33), .Y(
        n983) );
  OAI2BB2X1 U1995 ( .B0(n2225), .B1(n33), .A0N(\regs[28][2] ), .A1N(n33), .Y(
        n984) );
  OAI2BB2X1 U1996 ( .B0(n6), .B1(n33), .A0N(\regs[28][3] ), .A1N(n33), .Y(n985) );
  OAI2BB2X1 U1997 ( .B0(n7), .B1(n33), .A0N(\regs[28][4] ), .A1N(n33), .Y(n986) );
  OAI2BB2X1 U1998 ( .B0(n8), .B1(n33), .A0N(\regs[28][5] ), .A1N(n33), .Y(n987) );
  OAI2BB2X1 U1999 ( .B0(n9), .B1(n33), .A0N(\regs[28][6] ), .A1N(n33), .Y(n988) );
  OAI2BB2X1 U2000 ( .B0(n2221), .B1(n33), .A0N(\regs[28][13] ), .A1N(n33), .Y(
        n995) );
  OAI2BB2X1 U2001 ( .B0(n2218), .B1(n33), .A0N(\regs[28][16] ), .A1N(n33), .Y(
        n998) );
  OAI2BB2X1 U2002 ( .B0(n2217), .B1(n33), .A0N(\regs[28][17] ), .A1N(n33), .Y(
        n999) );
  OAI2BB2X1 U2003 ( .B0(n2216), .B1(n33), .A0N(\regs[28][18] ), .A1N(n33), .Y(
        n1000) );
  OAI2BB2X1 U2004 ( .B0(n2215), .B1(n33), .A0N(\regs[28][19] ), .A1N(n33), .Y(
        n1001) );
  OAI2BB2X1 U2005 ( .B0(n2214), .B1(n33), .A0N(\regs[28][20] ), .A1N(n33), .Y(
        n1002) );
  OAI2BB2X1 U2006 ( .B0(n2213), .B1(n33), .A0N(\regs[28][21] ), .A1N(n33), .Y(
        n1003) );
  OAI2BB2X1 U2007 ( .B0(n2212), .B1(n33), .A0N(\regs[28][22] ), .A1N(n33), .Y(
        n1004) );
  OAI2BB2X1 U2008 ( .B0(n2211), .B1(n33), .A0N(\regs[28][23] ), .A1N(n33), .Y(
        n1005) );
  OAI2BB2X1 U2009 ( .B0(n2210), .B1(n33), .A0N(\regs[28][24] ), .A1N(n33), .Y(
        n1006) );
  OAI2BB2X1 U2010 ( .B0(n2209), .B1(n33), .A0N(\regs[28][25] ), .A1N(n33), .Y(
        n1007) );
  OAI2BB2X1 U2011 ( .B0(n2208), .B1(n33), .A0N(\regs[28][26] ), .A1N(n33), .Y(
        n1008) );
  OAI2BB2X1 U2012 ( .B0(n2207), .B1(n33), .A0N(\regs[28][27] ), .A1N(n33), .Y(
        n1009) );
  OAI2BB2X1 U2013 ( .B0(n2206), .B1(n33), .A0N(\regs[28][28] ), .A1N(n33), .Y(
        n1010) );
  OAI2BB2X1 U2014 ( .B0(n2205), .B1(n33), .A0N(\regs[28][29] ), .A1N(n33), .Y(
        n1011) );
  OAI2BB2X1 U2015 ( .B0(n2204), .B1(n33), .A0N(\regs[28][30] ), .A1N(n33), .Y(
        n1012) );
  OAI2BB2X1 U2016 ( .B0(n34), .B1(n33), .A0N(\regs[28][31] ), .A1N(n33), .Y(
        n1013) );
  OAI2BB2X1 U2017 ( .B0(n2227), .B1(n37), .A0N(\regs[29][0] ), .A1N(n37), .Y(
        n1014) );
  OAI2BB2X1 U2018 ( .B0(n2226), .B1(n37), .A0N(\regs[29][1] ), .A1N(n37), .Y(
        n1015) );
  OAI2BB2X1 U2019 ( .B0(n2225), .B1(n37), .A0N(\regs[29][2] ), .A1N(n37), .Y(
        n1016) );
  OAI2BB2X1 U2020 ( .B0(n6), .B1(n37), .A0N(\regs[29][3] ), .A1N(n37), .Y(
        n1017) );
  OAI2BB2X1 U2021 ( .B0(n7), .B1(n37), .A0N(\regs[29][4] ), .A1N(n37), .Y(
        n1018) );
  OAI2BB2X1 U2022 ( .B0(n8), .B1(n37), .A0N(\regs[29][5] ), .A1N(n37), .Y(
        n1019) );
  OAI2BB2X1 U2023 ( .B0(n9), .B1(n37), .A0N(\regs[29][6] ), .A1N(n37), .Y(
        n1020) );
  OAI2BB2X1 U2024 ( .B0(n2221), .B1(n37), .A0N(\regs[29][13] ), .A1N(n37), .Y(
        n1027) );
  OAI2BB2X1 U2025 ( .B0(n2218), .B1(n37), .A0N(\regs[29][16] ), .A1N(n37), .Y(
        n1030) );
  OAI2BB2X1 U2026 ( .B0(n2217), .B1(n37), .A0N(\regs[29][17] ), .A1N(n37), .Y(
        n1031) );
  OAI2BB2X1 U2027 ( .B0(n2216), .B1(n37), .A0N(\regs[29][18] ), .A1N(n37), .Y(
        n1032) );
  OAI2BB2X1 U2028 ( .B0(n2215), .B1(n37), .A0N(\regs[29][19] ), .A1N(n37), .Y(
        n1033) );
  OAI2BB2X1 U2029 ( .B0(n2214), .B1(n37), .A0N(\regs[29][20] ), .A1N(n37), .Y(
        n1034) );
  OAI2BB2X1 U2030 ( .B0(n2213), .B1(n37), .A0N(\regs[29][21] ), .A1N(n37), .Y(
        n1035) );
  OAI2BB2X1 U2031 ( .B0(n2212), .B1(n37), .A0N(\regs[29][22] ), .A1N(n37), .Y(
        n1036) );
  OAI2BB2X1 U2032 ( .B0(n2211), .B1(n37), .A0N(\regs[29][23] ), .A1N(n37), .Y(
        n1037) );
  OAI2BB2X1 U2033 ( .B0(n2210), .B1(n37), .A0N(\regs[29][24] ), .A1N(n37), .Y(
        n1038) );
  OAI2BB2X1 U2034 ( .B0(n2209), .B1(n37), .A0N(\regs[29][25] ), .A1N(n37), .Y(
        n1039) );
  OAI2BB2X1 U2035 ( .B0(n2208), .B1(n37), .A0N(\regs[29][26] ), .A1N(n37), .Y(
        n1040) );
  OAI2BB2X1 U2036 ( .B0(n2207), .B1(n37), .A0N(\regs[29][27] ), .A1N(n37), .Y(
        n1041) );
  OAI2BB2X1 U2037 ( .B0(n2206), .B1(n37), .A0N(\regs[29][28] ), .A1N(n37), .Y(
        n1042) );
  OAI2BB2X1 U2038 ( .B0(n2205), .B1(n37), .A0N(\regs[29][29] ), .A1N(n37), .Y(
        n1043) );
  OAI2BB2X1 U2039 ( .B0(n2204), .B1(n37), .A0N(\regs[29][30] ), .A1N(n37), .Y(
        n1044) );
  OAI2BB2X1 U2040 ( .B0(n34), .B1(n37), .A0N(\regs[29][31] ), .A1N(n37), .Y(
        n1045) );
  OAI2BB2X1 U2041 ( .B0(n2227), .B1(n39), .A0N(\regs[30][0] ), .A1N(n39), .Y(
        n1046) );
  OAI2BB2X1 U2042 ( .B0(n2226), .B1(n39), .A0N(\regs[30][1] ), .A1N(n39), .Y(
        n1047) );
  OAI2BB2X1 U2043 ( .B0(n2225), .B1(n39), .A0N(\regs[30][2] ), .A1N(n39), .Y(
        n1048) );
  OAI2BB2X1 U2044 ( .B0(n6), .B1(n39), .A0N(\regs[30][3] ), .A1N(n39), .Y(
        n1049) );
  OAI2BB2X1 U2045 ( .B0(n7), .B1(n39), .A0N(\regs[30][4] ), .A1N(n39), .Y(
        n1050) );
  OAI2BB2X1 U2046 ( .B0(n8), .B1(n39), .A0N(\regs[30][5] ), .A1N(n39), .Y(
        n1051) );
  OAI2BB2X1 U2047 ( .B0(n9), .B1(n39), .A0N(\regs[30][6] ), .A1N(n39), .Y(
        n1052) );
  OAI2BB2X1 U2048 ( .B0(n2221), .B1(n39), .A0N(\regs[30][13] ), .A1N(n39), .Y(
        n1059) );
  OAI2BB2X1 U2049 ( .B0(n2218), .B1(n39), .A0N(\regs[30][16] ), .A1N(n39), .Y(
        n1062) );
  OAI2BB2X1 U2050 ( .B0(n2217), .B1(n39), .A0N(\regs[30][17] ), .A1N(n39), .Y(
        n1063) );
  OAI2BB2X1 U2051 ( .B0(n2216), .B1(n39), .A0N(\regs[30][18] ), .A1N(n39), .Y(
        n1064) );
  OAI2BB2X1 U2052 ( .B0(n2215), .B1(n39), .A0N(\regs[30][19] ), .A1N(n39), .Y(
        n1065) );
  OAI2BB2X1 U2053 ( .B0(n2214), .B1(n39), .A0N(\regs[30][20] ), .A1N(n39), .Y(
        n1066) );
  OAI2BB2X1 U2054 ( .B0(n2213), .B1(n39), .A0N(\regs[30][21] ), .A1N(n39), .Y(
        n1067) );
  OAI2BB2X1 U2055 ( .B0(n2212), .B1(n39), .A0N(\regs[30][22] ), .A1N(n39), .Y(
        n1068) );
  OAI2BB2X1 U2056 ( .B0(n2211), .B1(n39), .A0N(\regs[30][23] ), .A1N(n39), .Y(
        n1069) );
  OAI2BB2X1 U2057 ( .B0(n2210), .B1(n39), .A0N(\regs[30][24] ), .A1N(n39), .Y(
        n1070) );
  OAI2BB2X1 U2058 ( .B0(n2209), .B1(n39), .A0N(\regs[30][25] ), .A1N(n39), .Y(
        n1071) );
  OAI2BB2X1 U2059 ( .B0(n2208), .B1(n39), .A0N(\regs[30][26] ), .A1N(n39), .Y(
        n1072) );
  OAI2BB2X1 U2060 ( .B0(n2207), .B1(n39), .A0N(\regs[30][27] ), .A1N(n39), .Y(
        n1073) );
  OAI2BB2X1 U2061 ( .B0(n2206), .B1(n39), .A0N(\regs[30][28] ), .A1N(n39), .Y(
        n1074) );
  OAI2BB2X1 U2062 ( .B0(n2205), .B1(n39), .A0N(\regs[30][29] ), .A1N(n39), .Y(
        n1075) );
  OAI2BB2X1 U2063 ( .B0(n2204), .B1(n39), .A0N(\regs[30][30] ), .A1N(n39), .Y(
        n1076) );
  OAI2BB2X1 U2064 ( .B0(n34), .B1(n39), .A0N(\regs[30][31] ), .A1N(n39), .Y(
        n1077) );
  OAI2BB2X1 U2065 ( .B0(n2227), .B1(n41), .A0N(\regs[31][0] ), .A1N(n41), .Y(
        n1078) );
  OAI2BB2X1 U2066 ( .B0(n2226), .B1(n41), .A0N(\regs[31][1] ), .A1N(n41), .Y(
        n1079) );
  OAI2BB2X1 U2067 ( .B0(n2225), .B1(n41), .A0N(\regs[31][2] ), .A1N(n41), .Y(
        n1080) );
  OAI2BB2X1 U2068 ( .B0(n6), .B1(n41), .A0N(\regs[31][3] ), .A1N(n41), .Y(
        n1081) );
  OAI2BB2X1 U2069 ( .B0(n7), .B1(n41), .A0N(\regs[31][4] ), .A1N(n41), .Y(
        n1082) );
  OAI2BB2X1 U2070 ( .B0(n8), .B1(n41), .A0N(\regs[31][5] ), .A1N(n41), .Y(
        n1083) );
  OAI2BB2X1 U2071 ( .B0(n9), .B1(n41), .A0N(\regs[31][6] ), .A1N(n41), .Y(
        n1084) );
  OAI2BB2X1 U2072 ( .B0(n2221), .B1(n41), .A0N(\regs[31][13] ), .A1N(n41), .Y(
        n1091) );
  OAI2BB2X1 U2073 ( .B0(n2218), .B1(n41), .A0N(\regs[31][16] ), .A1N(n41), .Y(
        n1094) );
  OAI2BB2X1 U2074 ( .B0(n2217), .B1(n41), .A0N(\regs[31][17] ), .A1N(n41), .Y(
        n1095) );
  OAI2BB2X1 U2075 ( .B0(n2216), .B1(n41), .A0N(\regs[31][18] ), .A1N(n41), .Y(
        n1096) );
  OAI2BB2X1 U2076 ( .B0(n2215), .B1(n41), .A0N(\regs[31][19] ), .A1N(n41), .Y(
        n1097) );
  OAI2BB2X1 U2077 ( .B0(n2214), .B1(n41), .A0N(\regs[31][20] ), .A1N(n41), .Y(
        n1098) );
  OAI2BB2X1 U2078 ( .B0(n2213), .B1(n41), .A0N(\regs[31][21] ), .A1N(n41), .Y(
        n1099) );
  OAI2BB2X1 U2079 ( .B0(n2212), .B1(n41), .A0N(\regs[31][22] ), .A1N(n41), .Y(
        n1100) );
  OAI2BB2X1 U2080 ( .B0(n2211), .B1(n41), .A0N(\regs[31][23] ), .A1N(n41), .Y(
        n1101) );
  OAI2BB2X1 U2081 ( .B0(n2210), .B1(n41), .A0N(\regs[31][24] ), .A1N(n41), .Y(
        n1102) );
  OAI2BB2X1 U2082 ( .B0(n2209), .B1(n41), .A0N(\regs[31][25] ), .A1N(n41), .Y(
        n1103) );
  OAI2BB2X1 U2083 ( .B0(n2208), .B1(n41), .A0N(\regs[31][26] ), .A1N(n41), .Y(
        n1104) );
  OAI2BB2X1 U2084 ( .B0(n2207), .B1(n41), .A0N(\regs[31][27] ), .A1N(n41), .Y(
        n1105) );
  OAI2BB2X1 U2085 ( .B0(n2206), .B1(n41), .A0N(\regs[31][28] ), .A1N(n41), .Y(
        n1106) );
  OAI2BB2X1 U2086 ( .B0(n2205), .B1(n41), .A0N(\regs[31][29] ), .A1N(n41), .Y(
        n1107) );
  OAI2BB2X1 U2087 ( .B0(n2204), .B1(n41), .A0N(\regs[31][30] ), .A1N(n41), .Y(
        n1108) );
  OAI2BB2X1 U2088 ( .B0(n34), .B1(n41), .A0N(\regs[31][31] ), .A1N(n41), .Y(
        n1109) );
  OAI2BB2X1 U2089 ( .B0(n2), .B1(n2227), .A0N(\regs[0][0] ), .A1N(n2), .Y(n86)
         );
  OAI2BB2X1 U2090 ( .B0(n2), .B1(n2226), .A0N(\regs[0][1] ), .A1N(n2), .Y(n87)
         );
  OAI2BB2X1 U2091 ( .B0(n2), .B1(n2225), .A0N(\regs[0][2] ), .A1N(n2), .Y(n88)
         );
  OAI2BB2X1 U2092 ( .B0(n2), .B1(n6), .A0N(\regs[0][3] ), .A1N(n2), .Y(n89) );
  OAI2BB2X1 U2093 ( .B0(n2), .B1(n7), .A0N(\regs[0][4] ), .A1N(n2), .Y(n90) );
  OAI2BB2X1 U2094 ( .B0(n2), .B1(n8), .A0N(\regs[0][5] ), .A1N(n2), .Y(n91) );
  OAI2BB2X1 U2095 ( .B0(n2), .B1(n9), .A0N(\regs[0][6] ), .A1N(n2), .Y(n92) );
  OAI2BB2X1 U2096 ( .B0(n2), .B1(n10), .A0N(\regs[0][7] ), .A1N(n2), .Y(n93)
         );
  OAI2BB2X1 U2097 ( .B0(n2), .B1(n11), .A0N(\regs[0][8] ), .A1N(n2), .Y(n94)
         );
  OAI2BB2X1 U2098 ( .B0(n2), .B1(n12), .A0N(\regs[0][9] ), .A1N(n2), .Y(n95)
         );
  OAI2BB2X1 U2099 ( .B0(n2), .B1(n2224), .A0N(\regs[0][10] ), .A1N(n2), .Y(n96) );
  OAI2BB2X1 U2100 ( .B0(n2), .B1(n2223), .A0N(\regs[0][11] ), .A1N(n2), .Y(n97) );
  OAI2BB2X1 U2101 ( .B0(n2), .B1(n2222), .A0N(\regs[0][12] ), .A1N(n2), .Y(n98) );
  OAI2BB2X1 U2102 ( .B0(n2), .B1(n2221), .A0N(\regs[0][13] ), .A1N(n2), .Y(n99) );
  OAI2BB2X1 U2103 ( .B0(n2), .B1(n2220), .A0N(\regs[0][14] ), .A1N(n2), .Y(
        n100) );
  OAI2BB2X1 U2104 ( .B0(n2), .B1(n2219), .A0N(\regs[0][15] ), .A1N(n2), .Y(
        n101) );
  OAI2BB2X1 U2105 ( .B0(n2), .B1(n2218), .A0N(\regs[0][16] ), .A1N(n2), .Y(
        n102) );
  OAI2BB2X1 U2106 ( .B0(n2), .B1(n2217), .A0N(\regs[0][17] ), .A1N(n2), .Y(
        n103) );
  OAI2BB2X1 U2107 ( .B0(n2), .B1(n2216), .A0N(\regs[0][18] ), .A1N(n2), .Y(
        n104) );
  OAI2BB2X1 U2108 ( .B0(n2), .B1(n2215), .A0N(\regs[0][19] ), .A1N(n2), .Y(
        n105) );
  OAI2BB2X1 U2109 ( .B0(n2), .B1(n2214), .A0N(\regs[0][20] ), .A1N(n2), .Y(
        n106) );
  OAI2BB2X1 U2110 ( .B0(n2), .B1(n2213), .A0N(\regs[0][21] ), .A1N(n2), .Y(
        n107) );
  OAI2BB2X1 U2111 ( .B0(n2), .B1(n2212), .A0N(\regs[0][22] ), .A1N(n2), .Y(
        n108) );
  OAI2BB2X1 U2112 ( .B0(n2), .B1(n2211), .A0N(\regs[0][23] ), .A1N(n2), .Y(
        n109) );
  OAI2BB2X1 U2113 ( .B0(n2), .B1(n2210), .A0N(\regs[0][24] ), .A1N(n2), .Y(
        n110) );
  OAI2BB2X1 U2114 ( .B0(n2), .B1(n2209), .A0N(\regs[0][25] ), .A1N(n2), .Y(
        n111) );
  OAI2BB2X1 U2115 ( .B0(n2), .B1(n2208), .A0N(\regs[0][26] ), .A1N(n2), .Y(
        n112) );
  OAI2BB2X1 U2116 ( .B0(n2), .B1(n2207), .A0N(\regs[0][27] ), .A1N(n2), .Y(
        n113) );
  OAI2BB2X1 U2117 ( .B0(n2), .B1(n2206), .A0N(\regs[0][28] ), .A1N(n2), .Y(
        n114) );
  OAI2BB2X1 U2118 ( .B0(n2), .B1(n2205), .A0N(\regs[0][29] ), .A1N(n2), .Y(
        n115) );
  OAI2BB2X1 U2119 ( .B0(n2), .B1(n2204), .A0N(\regs[0][30] ), .A1N(n2), .Y(
        n116) );
  OAI2BB2X1 U2120 ( .B0(n2), .B1(n34), .A0N(\regs[0][31] ), .A1N(n2), .Y(n117)
         );
  MX4X1 U2121 ( .A(n1467), .B(n1465), .C(n1466), .D(n1464), .S0(N20), .S1(N19), 
        .Y(n1468) );
  MX4X1 U2122 ( .A(\regs[0][0] ), .B(\regs[1][0] ), .C(\regs[2][0] ), .D(
        \regs[3][0] ), .S0(n1809), .S1(n1786), .Y(n1467) );
  MX4X1 U2123 ( .A(\regs[8][0] ), .B(\regs[9][0] ), .C(\regs[10][0] ), .D(
        \regs[11][0] ), .S0(n1809), .S1(n1786), .Y(n1465) );
  MX4X1 U2124 ( .A(\regs[4][0] ), .B(\regs[5][0] ), .C(\regs[6][0] ), .D(
        \regs[7][0] ), .S0(n1809), .S1(n1786), .Y(n1466) );
  MX4X1 U2125 ( .A(\regs[20][0] ), .B(\regs[21][0] ), .C(\regs[22][0] ), .D(
        \regs[23][0] ), .S0(n1808), .S1(n1798), .Y(n1461) );
  MX4X1 U2126 ( .A(\regs[4][1] ), .B(\regs[5][1] ), .C(\regs[6][1] ), .D(
        \regs[7][1] ), .S0(n1809), .S1(n1786), .Y(n1476) );
  MX4X1 U2127 ( .A(\regs[4][2] ), .B(\regs[5][2] ), .C(\regs[6][2] ), .D(
        \regs[7][2] ), .S0(n1810), .S1(n1787), .Y(n1486) );
  MX4X1 U2128 ( .A(\regs[4][3] ), .B(\regs[5][3] ), .C(\regs[6][3] ), .D(
        \regs[7][3] ), .S0(n1811), .S1(n1788), .Y(n1496) );
  MX4X1 U2129 ( .A(\regs[4][4] ), .B(\regs[5][4] ), .C(\regs[6][4] ), .D(
        \regs[7][4] ), .S0(n1811), .S1(n1788), .Y(n1506) );
  MX4X1 U2130 ( .A(\regs[4][5] ), .B(\regs[5][5] ), .C(\regs[6][5] ), .D(
        \regs[7][5] ), .S0(n1812), .S1(n1789), .Y(n1516) );
  MX4X1 U2131 ( .A(\regs[4][6] ), .B(\regs[5][6] ), .C(\regs[6][6] ), .D(
        \regs[7][6] ), .S0(n1813), .S1(n1790), .Y(n1526) );
  MX4X1 U2132 ( .A(\regs[4][7] ), .B(\regs[5][7] ), .C(\regs[6][7] ), .D(
        \regs[7][7] ), .S0(n1813), .S1(n1790), .Y(n1536) );
  MX4X1 U2133 ( .A(\regs[4][8] ), .B(\regs[5][8] ), .C(\regs[6][8] ), .D(
        \regs[7][8] ), .S0(n1814), .S1(n1791), .Y(n1546) );
  MX4X1 U2134 ( .A(\regs[4][9] ), .B(\regs[5][9] ), .C(\regs[6][9] ), .D(
        \regs[7][9] ), .S0(n1815), .S1(n1792), .Y(n1556) );
  MX4X1 U2135 ( .A(\regs[4][10] ), .B(\regs[5][10] ), .C(\regs[6][10] ), .D(
        \regs[7][10] ), .S0(n1815), .S1(n1792), .Y(n1566) );
  MX4X1 U2136 ( .A(\regs[4][11] ), .B(\regs[5][11] ), .C(\regs[6][11] ), .D(
        \regs[7][11] ), .S0(n1816), .S1(n1793), .Y(n1576) );
  MX4X1 U2137 ( .A(\regs[4][12] ), .B(\regs[5][12] ), .C(\regs[6][12] ), .D(
        \regs[7][12] ), .S0(n1817), .S1(n1794), .Y(n1586) );
  MX4X1 U2138 ( .A(\regs[4][13] ), .B(\regs[5][13] ), .C(\regs[6][13] ), .D(
        \regs[7][13] ), .S0(n1817), .S1(n1794), .Y(n1596) );
  MX4X1 U2139 ( .A(\regs[4][14] ), .B(\regs[5][14] ), .C(\regs[6][14] ), .D(
        \regs[7][14] ), .S0(n1818), .S1(n1795), .Y(n1606) );
  MX4X1 U2140 ( .A(\regs[4][15] ), .B(\regs[5][15] ), .C(\regs[6][15] ), .D(
        \regs[7][15] ), .S0(n1819), .S1(n1796), .Y(n1616) );
  MX4X1 U2141 ( .A(\regs[4][16] ), .B(\regs[5][16] ), .C(\regs[6][16] ), .D(
        \regs[7][16] ), .S0(n1819), .S1(n1796), .Y(n1626) );
  MX4X1 U2142 ( .A(\regs[4][17] ), .B(\regs[5][17] ), .C(\regs[6][17] ), .D(
        \regs[7][17] ), .S0(n1820), .S1(n1797), .Y(n1636) );
  MX4X1 U2143 ( .A(\regs[4][18] ), .B(\regs[5][18] ), .C(\regs[6][18] ), .D(
        \regs[7][18] ), .S0(n1821), .S1(n1798), .Y(n1646) );
  MX4X1 U2144 ( .A(\regs[4][19] ), .B(\regs[5][19] ), .C(\regs[6][19] ), .D(
        \regs[7][19] ), .S0(n1821), .S1(n1798), .Y(n1656) );
  MX4X1 U2145 ( .A(\regs[4][20] ), .B(\regs[5][20] ), .C(\regs[6][20] ), .D(
        \regs[7][20] ), .S0(n1822), .S1(n1799), .Y(n1666) );
  MX4X1 U2146 ( .A(\regs[4][21] ), .B(\regs[5][21] ), .C(\regs[6][21] ), .D(
        \regs[7][21] ), .S0(n1823), .S1(n1800), .Y(n1676) );
  MX4X1 U2147 ( .A(\regs[4][22] ), .B(\regs[5][22] ), .C(\regs[6][22] ), .D(
        \regs[7][22] ), .S0(n1823), .S1(n1800), .Y(n1686) );
  MX4X1 U2148 ( .A(\regs[4][23] ), .B(\regs[5][23] ), .C(\regs[6][23] ), .D(
        \regs[7][23] ), .S0(n1824), .S1(n1801), .Y(n1696) );
  MX4X1 U2149 ( .A(\regs[4][24] ), .B(\regs[5][24] ), .C(\regs[6][24] ), .D(
        \regs[7][24] ), .S0(n1825), .S1(n1802), .Y(n1706) );
  MX4X1 U2150 ( .A(\regs[4][25] ), .B(\regs[5][25] ), .C(\regs[6][25] ), .D(
        \regs[7][25] ), .S0(n1825), .S1(n1802), .Y(n1716) );
  MX4X1 U2151 ( .A(\regs[4][26] ), .B(\regs[5][26] ), .C(\regs[6][26] ), .D(
        \regs[7][26] ), .S0(n1826), .S1(n1803), .Y(n1726) );
  MX4X1 U2152 ( .A(\regs[4][27] ), .B(\regs[5][27] ), .C(\regs[6][27] ), .D(
        \regs[7][27] ), .S0(n1827), .S1(n1804), .Y(n1736) );
  MX4X1 U2153 ( .A(\regs[4][28] ), .B(\regs[5][28] ), .C(\regs[6][28] ), .D(
        \regs[7][28] ), .S0(n1827), .S1(n1804), .Y(n1746) );
  MX4X1 U2154 ( .A(\regs[4][29] ), .B(\regs[5][29] ), .C(\regs[6][29] ), .D(
        \regs[7][29] ), .S0(n1828), .S1(n1805), .Y(n1756) );
  MX4X1 U2155 ( .A(\regs[4][30] ), .B(\regs[5][30] ), .C(\regs[6][30] ), .D(
        \regs[7][30] ), .S0(n1829), .S1(n1806), .Y(n1766) );
  MX4X1 U2156 ( .A(\regs[4][31] ), .B(\regs[5][31] ), .C(\regs[6][31] ), .D(
        \regs[7][31] ), .S0(n1829), .S1(n1806), .Y(n1776) );
  MX4X1 U2157 ( .A(\regs[16][0] ), .B(\regs[17][0] ), .C(\regs[18][0] ), .D(
        \regs[19][0] ), .S0(n1808), .S1(n1786), .Y(n1462) );
  MX4X1 U2158 ( .A(\regs[0][1] ), .B(\regs[1][1] ), .C(\regs[2][1] ), .D(
        \regs[3][1] ), .S0(n1809), .S1(n1786), .Y(n1477) );
  MX4X1 U2159 ( .A(\regs[0][2] ), .B(\regs[1][2] ), .C(\regs[2][2] ), .D(
        \regs[3][2] ), .S0(n1810), .S1(n1787), .Y(n1487) );
  MX4X1 U2160 ( .A(\regs[0][3] ), .B(\regs[1][3] ), .C(\regs[2][3] ), .D(
        \regs[3][3] ), .S0(n1811), .S1(n1788), .Y(n1497) );
  MX4X1 U2161 ( .A(\regs[0][4] ), .B(\regs[1][4] ), .C(\regs[2][4] ), .D(
        \regs[3][4] ), .S0(n1811), .S1(n1788), .Y(n1507) );
  MX4X1 U2162 ( .A(\regs[0][5] ), .B(\regs[1][5] ), .C(\regs[2][5] ), .D(
        \regs[3][5] ), .S0(n1812), .S1(n1789), .Y(n1517) );
  MX4X1 U2163 ( .A(\regs[0][6] ), .B(\regs[1][6] ), .C(\regs[2][6] ), .D(
        \regs[3][6] ), .S0(n1813), .S1(n1790), .Y(n1527) );
  MX4X1 U2164 ( .A(\regs[0][7] ), .B(\regs[1][7] ), .C(\regs[2][7] ), .D(
        \regs[3][7] ), .S0(n1813), .S1(n1790), .Y(n1537) );
  MX4X1 U2165 ( .A(\regs[0][8] ), .B(\regs[1][8] ), .C(\regs[2][8] ), .D(
        \regs[3][8] ), .S0(n1814), .S1(n1791), .Y(n1547) );
  MX4X1 U2166 ( .A(\regs[0][9] ), .B(\regs[1][9] ), .C(\regs[2][9] ), .D(
        \regs[3][9] ), .S0(n1815), .S1(n1792), .Y(n1557) );
  MX4X1 U2167 ( .A(\regs[0][10] ), .B(\regs[1][10] ), .C(\regs[2][10] ), .D(
        \regs[3][10] ), .S0(n1815), .S1(n1792), .Y(n1567) );
  MX4X1 U2168 ( .A(\regs[0][11] ), .B(\regs[1][11] ), .C(\regs[2][11] ), .D(
        \regs[3][11] ), .S0(n1816), .S1(n1793), .Y(n1577) );
  MX4X1 U2169 ( .A(\regs[0][12] ), .B(\regs[1][12] ), .C(\regs[2][12] ), .D(
        \regs[3][12] ), .S0(n1817), .S1(n1794), .Y(n1587) );
  MX4X1 U2170 ( .A(\regs[0][13] ), .B(\regs[1][13] ), .C(\regs[2][13] ), .D(
        \regs[3][13] ), .S0(n1817), .S1(n1794), .Y(n1597) );
  MX4X1 U2171 ( .A(\regs[0][14] ), .B(\regs[1][14] ), .C(\regs[2][14] ), .D(
        \regs[3][14] ), .S0(n1818), .S1(n1795), .Y(n1607) );
  MX4X1 U2172 ( .A(\regs[0][15] ), .B(\regs[1][15] ), .C(\regs[2][15] ), .D(
        \regs[3][15] ), .S0(n1819), .S1(n1796), .Y(n1617) );
  MX4X1 U2173 ( .A(\regs[0][16] ), .B(\regs[1][16] ), .C(\regs[2][16] ), .D(
        \regs[3][16] ), .S0(n1819), .S1(n1796), .Y(n1627) );
  MX4X1 U2174 ( .A(\regs[0][17] ), .B(\regs[1][17] ), .C(\regs[2][17] ), .D(
        \regs[3][17] ), .S0(n1820), .S1(n1797), .Y(n1637) );
  MX4X1 U2175 ( .A(\regs[0][18] ), .B(\regs[1][18] ), .C(\regs[2][18] ), .D(
        \regs[3][18] ), .S0(n1821), .S1(n1798), .Y(n1647) );
  MX4X1 U2176 ( .A(\regs[0][19] ), .B(\regs[1][19] ), .C(\regs[2][19] ), .D(
        \regs[3][19] ), .S0(n1821), .S1(n1798), .Y(n1657) );
  MX4X1 U2177 ( .A(\regs[0][20] ), .B(\regs[1][20] ), .C(\regs[2][20] ), .D(
        \regs[3][20] ), .S0(n1822), .S1(n1799), .Y(n1667) );
  MX4X1 U2178 ( .A(\regs[0][21] ), .B(\regs[1][21] ), .C(\regs[2][21] ), .D(
        \regs[3][21] ), .S0(n1823), .S1(n1800), .Y(n1677) );
  MX4X1 U2179 ( .A(\regs[0][22] ), .B(\regs[1][22] ), .C(\regs[2][22] ), .D(
        \regs[3][22] ), .S0(n1823), .S1(n1800), .Y(n1687) );
  MX4X1 U2180 ( .A(\regs[0][23] ), .B(\regs[1][23] ), .C(\regs[2][23] ), .D(
        \regs[3][23] ), .S0(n1824), .S1(n1801), .Y(n1697) );
  MX4X1 U2181 ( .A(\regs[0][24] ), .B(\regs[1][24] ), .C(\regs[2][24] ), .D(
        \regs[3][24] ), .S0(n1825), .S1(n1802), .Y(n1707) );
  MX4X1 U2182 ( .A(\regs[0][25] ), .B(\regs[1][25] ), .C(\regs[2][25] ), .D(
        \regs[3][25] ), .S0(n1825), .S1(n1802), .Y(n1717) );
  MX4X1 U2183 ( .A(\regs[0][26] ), .B(\regs[1][26] ), .C(\regs[2][26] ), .D(
        \regs[3][26] ), .S0(n1826), .S1(n1803), .Y(n1727) );
  MX4X1 U2184 ( .A(\regs[0][27] ), .B(\regs[1][27] ), .C(\regs[2][27] ), .D(
        \regs[3][27] ), .S0(n1827), .S1(n1804), .Y(n1737) );
  MX4X1 U2185 ( .A(\regs[0][28] ), .B(\regs[1][28] ), .C(\regs[2][28] ), .D(
        \regs[3][28] ), .S0(n1827), .S1(n1804), .Y(n1747) );
  MX4X1 U2186 ( .A(\regs[0][29] ), .B(\regs[1][29] ), .C(\regs[2][29] ), .D(
        \regs[3][29] ), .S0(n1828), .S1(n1805), .Y(n1757) );
  MX4X1 U2187 ( .A(\regs[0][30] ), .B(\regs[1][30] ), .C(\regs[2][30] ), .D(
        \regs[3][30] ), .S0(n1829), .S1(n1806), .Y(n1767) );
  MX4X1 U2188 ( .A(\regs[0][31] ), .B(\regs[1][31] ), .C(\regs[2][31] ), .D(
        \regs[3][31] ), .S0(n1829), .S1(n1806), .Y(n1777) );
  MX4X1 U2189 ( .A(\regs[12][0] ), .B(\regs[13][0] ), .C(\regs[14][0] ), .D(
        \regs[15][0] ), .S0(n1809), .S1(n1786), .Y(n1464) );
  MX4X1 U2190 ( .A(\regs[28][0] ), .B(\regs[29][0] ), .C(\regs[30][0] ), .D(
        \regs[31][0] ), .S0(n1808), .S1(n1796), .Y(n1459) );
  MX4X1 U2191 ( .A(\regs[28][1] ), .B(\regs[29][1] ), .C(\regs[30][1] ), .D(
        \regs[31][1] ), .S0(n1809), .S1(n1786), .Y(n1469) );
  MX4X1 U2192 ( .A(\regs[12][1] ), .B(\regs[13][1] ), .C(\regs[14][1] ), .D(
        \regs[15][1] ), .S0(n1809), .S1(n1786), .Y(n1474) );
  MX4X1 U2193 ( .A(\regs[28][2] ), .B(\regs[29][2] ), .C(\regs[30][2] ), .D(
        \regs[31][2] ), .S0(n1810), .S1(n1787), .Y(n1479) );
  MX4X1 U2194 ( .A(\regs[12][2] ), .B(\regs[13][2] ), .C(\regs[14][2] ), .D(
        \regs[15][2] ), .S0(n1810), .S1(n1787), .Y(n1484) );
  MX4X1 U2195 ( .A(\regs[28][3] ), .B(\regs[29][3] ), .C(\regs[30][3] ), .D(
        \regs[31][3] ), .S0(n1810), .S1(n1787), .Y(n1489) );
  MX4X1 U2196 ( .A(\regs[12][3] ), .B(\regs[13][3] ), .C(\regs[14][3] ), .D(
        \regs[15][3] ), .S0(n1811), .S1(n1788), .Y(n1494) );
  MX4X1 U2197 ( .A(\regs[28][4] ), .B(\regs[29][4] ), .C(\regs[30][4] ), .D(
        \regs[31][4] ), .S0(n1811), .S1(n1788), .Y(n1499) );
  MX4X1 U2198 ( .A(\regs[12][4] ), .B(\regs[13][4] ), .C(\regs[14][4] ), .D(
        \regs[15][4] ), .S0(n1811), .S1(n1788), .Y(n1504) );
  MX4X1 U2199 ( .A(\regs[28][5] ), .B(\regs[29][5] ), .C(\regs[30][5] ), .D(
        \regs[31][5] ), .S0(n1812), .S1(n1789), .Y(n1509) );
  MX4X1 U2200 ( .A(\regs[12][5] ), .B(\regs[13][5] ), .C(\regs[14][5] ), .D(
        \regs[15][5] ), .S0(n1812), .S1(n1789), .Y(n1514) );
  MX4X1 U2201 ( .A(\regs[28][6] ), .B(\regs[29][6] ), .C(\regs[30][6] ), .D(
        \regs[31][6] ), .S0(n1812), .S1(n1789), .Y(n1519) );
  MX4X1 U2202 ( .A(\regs[12][6] ), .B(\regs[13][6] ), .C(\regs[14][6] ), .D(
        \regs[15][6] ), .S0(n1813), .S1(n1790), .Y(n1524) );
  MX4X1 U2203 ( .A(\regs[28][7] ), .B(\regs[29][7] ), .C(\regs[30][7] ), .D(
        \regs[31][7] ), .S0(n1813), .S1(n1790), .Y(n1529) );
  MX4X1 U2204 ( .A(\regs[12][7] ), .B(\regs[13][7] ), .C(\regs[14][7] ), .D(
        \regs[15][7] ), .S0(n1813), .S1(n1790), .Y(n1534) );
  MX4X1 U2205 ( .A(\regs[28][8] ), .B(\regs[29][8] ), .C(\regs[30][8] ), .D(
        \regs[31][8] ), .S0(n1814), .S1(n1791), .Y(n1539) );
  MX4X1 U2206 ( .A(\regs[12][8] ), .B(\regs[13][8] ), .C(\regs[14][8] ), .D(
        \regs[15][8] ), .S0(n1814), .S1(n1791), .Y(n1544) );
  MX4X1 U2207 ( .A(\regs[28][9] ), .B(\regs[29][9] ), .C(\regs[30][9] ), .D(
        \regs[31][9] ), .S0(n1814), .S1(n1791), .Y(n1549) );
  MX4X1 U2208 ( .A(\regs[12][9] ), .B(\regs[13][9] ), .C(\regs[14][9] ), .D(
        \regs[15][9] ), .S0(n1815), .S1(n1792), .Y(n1554) );
  MX4X1 U2209 ( .A(\regs[28][10] ), .B(\regs[29][10] ), .C(\regs[30][10] ), 
        .D(\regs[31][10] ), .S0(n1815), .S1(n1792), .Y(n1559) );
  MX4X1 U2210 ( .A(\regs[12][10] ), .B(\regs[13][10] ), .C(\regs[14][10] ), 
        .D(\regs[15][10] ), .S0(n1815), .S1(n1792), .Y(n1564) );
  MX4X1 U2211 ( .A(\regs[28][11] ), .B(\regs[29][11] ), .C(\regs[30][11] ), 
        .D(\regs[31][11] ), .S0(n1816), .S1(n1793), .Y(n1569) );
  MX4X1 U2212 ( .A(\regs[12][11] ), .B(\regs[13][11] ), .C(\regs[14][11] ), 
        .D(\regs[15][11] ), .S0(n1816), .S1(n1793), .Y(n1574) );
  MX4X1 U2213 ( .A(\regs[28][12] ), .B(\regs[29][12] ), .C(\regs[30][12] ), 
        .D(\regs[31][12] ), .S0(n1816), .S1(n1793), .Y(n1579) );
  MX4X1 U2214 ( .A(\regs[12][12] ), .B(\regs[13][12] ), .C(\regs[14][12] ), 
        .D(\regs[15][12] ), .S0(n1817), .S1(n1794), .Y(n1584) );
  MX4X1 U2215 ( .A(\regs[28][13] ), .B(\regs[29][13] ), .C(\regs[30][13] ), 
        .D(\regs[31][13] ), .S0(n1817), .S1(n1794), .Y(n1589) );
  MX4X1 U2216 ( .A(\regs[12][13] ), .B(\regs[13][13] ), .C(\regs[14][13] ), 
        .D(\regs[15][13] ), .S0(n1817), .S1(n1794), .Y(n1594) );
  MX4X1 U2217 ( .A(\regs[28][14] ), .B(\regs[29][14] ), .C(\regs[30][14] ), 
        .D(\regs[31][14] ), .S0(n1818), .S1(n1795), .Y(n1599) );
  MX4X1 U2218 ( .A(\regs[12][14] ), .B(\regs[13][14] ), .C(\regs[14][14] ), 
        .D(\regs[15][14] ), .S0(n1818), .S1(n1795), .Y(n1604) );
  MX4X1 U2219 ( .A(\regs[28][15] ), .B(\regs[29][15] ), .C(\regs[30][15] ), 
        .D(\regs[31][15] ), .S0(n1818), .S1(n1795), .Y(n1609) );
  MX4X1 U2220 ( .A(\regs[12][15] ), .B(\regs[13][15] ), .C(\regs[14][15] ), 
        .D(\regs[15][15] ), .S0(n1819), .S1(n1796), .Y(n1614) );
  MX4X1 U2221 ( .A(\regs[28][16] ), .B(\regs[29][16] ), .C(\regs[30][16] ), 
        .D(\regs[31][16] ), .S0(n1819), .S1(n1796), .Y(n1619) );
  MX4X1 U2222 ( .A(\regs[12][16] ), .B(\regs[13][16] ), .C(\regs[14][16] ), 
        .D(\regs[15][16] ), .S0(n1819), .S1(n1796), .Y(n1624) );
  MX4X1 U2223 ( .A(\regs[28][17] ), .B(\regs[29][17] ), .C(\regs[30][17] ), 
        .D(\regs[31][17] ), .S0(n1820), .S1(n1797), .Y(n1629) );
  MX4X1 U2224 ( .A(\regs[12][17] ), .B(\regs[13][17] ), .C(\regs[14][17] ), 
        .D(\regs[15][17] ), .S0(n1820), .S1(n1797), .Y(n1634) );
  MX4X1 U2225 ( .A(\regs[28][18] ), .B(\regs[29][18] ), .C(\regs[30][18] ), 
        .D(\regs[31][18] ), .S0(n1820), .S1(n1797), .Y(n1639) );
  MX4X1 U2226 ( .A(\regs[12][18] ), .B(\regs[13][18] ), .C(\regs[14][18] ), 
        .D(\regs[15][18] ), .S0(n1821), .S1(n1798), .Y(n1644) );
  MX4X1 U2227 ( .A(\regs[28][19] ), .B(\regs[29][19] ), .C(\regs[30][19] ), 
        .D(\regs[31][19] ), .S0(n1821), .S1(n1798), .Y(n1649) );
  MX4X1 U2228 ( .A(\regs[12][19] ), .B(\regs[13][19] ), .C(\regs[14][19] ), 
        .D(\regs[15][19] ), .S0(n1821), .S1(n1798), .Y(n1654) );
  MX4X1 U2229 ( .A(\regs[28][20] ), .B(\regs[29][20] ), .C(\regs[30][20] ), 
        .D(\regs[31][20] ), .S0(n1822), .S1(n1799), .Y(n1659) );
  MX4X1 U2230 ( .A(\regs[12][20] ), .B(\regs[13][20] ), .C(\regs[14][20] ), 
        .D(\regs[15][20] ), .S0(n1822), .S1(n1799), .Y(n1664) );
  MX4X1 U2231 ( .A(\regs[28][21] ), .B(\regs[29][21] ), .C(\regs[30][21] ), 
        .D(\regs[31][21] ), .S0(n1822), .S1(n1799), .Y(n1669) );
  MX4X1 U2232 ( .A(\regs[12][21] ), .B(\regs[13][21] ), .C(\regs[14][21] ), 
        .D(\regs[15][21] ), .S0(n1823), .S1(n1800), .Y(n1674) );
  MX4X1 U2233 ( .A(\regs[28][22] ), .B(\regs[29][22] ), .C(\regs[30][22] ), 
        .D(\regs[31][22] ), .S0(n1823), .S1(n1800), .Y(n1679) );
  MX4X1 U2234 ( .A(\regs[12][22] ), .B(\regs[13][22] ), .C(\regs[14][22] ), 
        .D(\regs[15][22] ), .S0(n1823), .S1(n1800), .Y(n1684) );
  MX4X1 U2235 ( .A(\regs[28][23] ), .B(\regs[29][23] ), .C(\regs[30][23] ), 
        .D(\regs[31][23] ), .S0(n1824), .S1(n1801), .Y(n1689) );
  MX4X1 U2236 ( .A(\regs[12][23] ), .B(\regs[13][23] ), .C(\regs[14][23] ), 
        .D(\regs[15][23] ), .S0(n1824), .S1(n1801), .Y(n1694) );
  MX4X1 U2237 ( .A(\regs[28][24] ), .B(\regs[29][24] ), .C(\regs[30][24] ), 
        .D(\regs[31][24] ), .S0(n1824), .S1(n1801), .Y(n1699) );
  MX4X1 U2238 ( .A(\regs[12][24] ), .B(\regs[13][24] ), .C(\regs[14][24] ), 
        .D(\regs[15][24] ), .S0(n1825), .S1(n1802), .Y(n1704) );
  MX4X1 U2239 ( .A(\regs[28][25] ), .B(\regs[29][25] ), .C(\regs[30][25] ), 
        .D(\regs[31][25] ), .S0(n1825), .S1(n1802), .Y(n1709) );
  MX4X1 U2240 ( .A(\regs[12][25] ), .B(\regs[13][25] ), .C(\regs[14][25] ), 
        .D(\regs[15][25] ), .S0(n1825), .S1(n1802), .Y(n1714) );
  MX4X1 U2241 ( .A(\regs[28][26] ), .B(\regs[29][26] ), .C(\regs[30][26] ), 
        .D(\regs[31][26] ), .S0(n1826), .S1(n1803), .Y(n1719) );
  MX4X1 U2242 ( .A(\regs[12][26] ), .B(\regs[13][26] ), .C(\regs[14][26] ), 
        .D(\regs[15][26] ), .S0(n1826), .S1(n1803), .Y(n1724) );
  MX4X1 U2243 ( .A(\regs[28][27] ), .B(\regs[29][27] ), .C(\regs[30][27] ), 
        .D(\regs[31][27] ), .S0(n1826), .S1(n1803), .Y(n1729) );
  MX4X1 U2244 ( .A(\regs[12][27] ), .B(\regs[13][27] ), .C(\regs[14][27] ), 
        .D(\regs[15][27] ), .S0(n1827), .S1(n1804), .Y(n1734) );
  MX4X1 U2245 ( .A(\regs[28][28] ), .B(\regs[29][28] ), .C(\regs[30][28] ), 
        .D(\regs[31][28] ), .S0(n1827), .S1(n1804), .Y(n1739) );
  MX4X1 U2246 ( .A(\regs[12][28] ), .B(\regs[13][28] ), .C(\regs[14][28] ), 
        .D(\regs[15][28] ), .S0(n1827), .S1(n1804), .Y(n1744) );
  MX4X1 U2247 ( .A(\regs[28][29] ), .B(\regs[29][29] ), .C(\regs[30][29] ), 
        .D(\regs[31][29] ), .S0(n1828), .S1(n1805), .Y(n1749) );
  MX4X1 U2248 ( .A(\regs[12][29] ), .B(\regs[13][29] ), .C(\regs[14][29] ), 
        .D(\regs[15][29] ), .S0(n1828), .S1(n1805), .Y(n1754) );
  MX4X1 U2249 ( .A(\regs[28][30] ), .B(\regs[29][30] ), .C(\regs[30][30] ), 
        .D(\regs[31][30] ), .S0(n1828), .S1(n1805), .Y(n1759) );
  MX4X1 U2250 ( .A(\regs[12][30] ), .B(\regs[13][30] ), .C(\regs[14][30] ), 
        .D(\regs[15][30] ), .S0(n1829), .S1(n1806), .Y(n1764) );
  MX4X1 U2251 ( .A(\regs[28][31] ), .B(\regs[29][31] ), .C(\regs[30][31] ), 
        .D(\regs[31][31] ), .S0(n1829), .S1(n1806), .Y(n1769) );
  MX4X1 U2252 ( .A(\regs[12][31] ), .B(\regs[13][31] ), .C(\regs[14][31] ), 
        .D(\regs[15][31] ), .S0(n1829), .S1(n1806), .Y(n1774) );
  MX4X1 U2253 ( .A(\regs[24][0] ), .B(\regs[25][0] ), .C(\regs[26][0] ), .D(
        \regs[27][0] ), .S0(n1808), .S1(n1795), .Y(n1460) );
  MX4X1 U2254 ( .A(\regs[8][1] ), .B(\regs[9][1] ), .C(\regs[10][1] ), .D(
        \regs[11][1] ), .S0(n1809), .S1(n1786), .Y(n1475) );
  MX4X1 U2255 ( .A(\regs[8][2] ), .B(\regs[9][2] ), .C(\regs[10][2] ), .D(
        \regs[11][2] ), .S0(n1810), .S1(n1787), .Y(n1485) );
  MX4X1 U2256 ( .A(\regs[8][3] ), .B(\regs[9][3] ), .C(\regs[10][3] ), .D(
        \regs[11][3] ), .S0(n1811), .S1(n1788), .Y(n1495) );
  MX4X1 U2257 ( .A(\regs[8][4] ), .B(\regs[9][4] ), .C(\regs[10][4] ), .D(
        \regs[11][4] ), .S0(n1811), .S1(n1788), .Y(n1505) );
  MX4X1 U2258 ( .A(\regs[8][5] ), .B(\regs[9][5] ), .C(\regs[10][5] ), .D(
        \regs[11][5] ), .S0(n1812), .S1(n1789), .Y(n1515) );
  MX4X1 U2259 ( .A(\regs[8][6] ), .B(\regs[9][6] ), .C(\regs[10][6] ), .D(
        \regs[11][6] ), .S0(n1813), .S1(n1790), .Y(n1525) );
  MX4X1 U2260 ( .A(\regs[8][7] ), .B(\regs[9][7] ), .C(\regs[10][7] ), .D(
        \regs[11][7] ), .S0(n1813), .S1(n1790), .Y(n1535) );
  MX4X1 U2261 ( .A(\regs[8][8] ), .B(\regs[9][8] ), .C(\regs[10][8] ), .D(
        \regs[11][8] ), .S0(n1814), .S1(n1791), .Y(n1545) );
  MX4X1 U2262 ( .A(\regs[8][9] ), .B(\regs[9][9] ), .C(\regs[10][9] ), .D(
        \regs[11][9] ), .S0(n1815), .S1(n1792), .Y(n1555) );
  MX4X1 U2263 ( .A(\regs[8][10] ), .B(\regs[9][10] ), .C(\regs[10][10] ), .D(
        \regs[11][10] ), .S0(n1815), .S1(n1792), .Y(n1565) );
  MX4X1 U2264 ( .A(\regs[8][11] ), .B(\regs[9][11] ), .C(\regs[10][11] ), .D(
        \regs[11][11] ), .S0(n1816), .S1(n1793), .Y(n1575) );
  MX4X1 U2265 ( .A(\regs[8][12] ), .B(\regs[9][12] ), .C(\regs[10][12] ), .D(
        \regs[11][12] ), .S0(n1817), .S1(n1794), .Y(n1585) );
  MX4X1 U2266 ( .A(\regs[8][13] ), .B(\regs[9][13] ), .C(\regs[10][13] ), .D(
        \regs[11][13] ), .S0(n1817), .S1(n1794), .Y(n1595) );
  MX4X1 U2267 ( .A(\regs[8][14] ), .B(\regs[9][14] ), .C(\regs[10][14] ), .D(
        \regs[11][14] ), .S0(n1818), .S1(n1795), .Y(n1605) );
  MX4X1 U2268 ( .A(\regs[8][15] ), .B(\regs[9][15] ), .C(\regs[10][15] ), .D(
        \regs[11][15] ), .S0(n1819), .S1(n1796), .Y(n1615) );
  MX4X1 U2269 ( .A(\regs[8][16] ), .B(\regs[9][16] ), .C(\regs[10][16] ), .D(
        \regs[11][16] ), .S0(n1819), .S1(n1796), .Y(n1625) );
  MX4X1 U2270 ( .A(\regs[8][17] ), .B(\regs[9][17] ), .C(\regs[10][17] ), .D(
        \regs[11][17] ), .S0(n1820), .S1(n1797), .Y(n1635) );
  MX4X1 U2271 ( .A(\regs[8][18] ), .B(\regs[9][18] ), .C(\regs[10][18] ), .D(
        \regs[11][18] ), .S0(n1821), .S1(n1798), .Y(n1645) );
  MX4X1 U2272 ( .A(\regs[8][19] ), .B(\regs[9][19] ), .C(\regs[10][19] ), .D(
        \regs[11][19] ), .S0(n1821), .S1(n1798), .Y(n1655) );
  MX4X1 U2273 ( .A(\regs[8][20] ), .B(\regs[9][20] ), .C(\regs[10][20] ), .D(
        \regs[11][20] ), .S0(n1822), .S1(n1799), .Y(n1665) );
  MX4X1 U2274 ( .A(\regs[8][21] ), .B(\regs[9][21] ), .C(\regs[10][21] ), .D(
        \regs[11][21] ), .S0(n1823), .S1(n1800), .Y(n1675) );
  MX4X1 U2275 ( .A(\regs[8][22] ), .B(\regs[9][22] ), .C(\regs[10][22] ), .D(
        \regs[11][22] ), .S0(n1823), .S1(n1800), .Y(n1685) );
  MX4X1 U2276 ( .A(\regs[8][23] ), .B(\regs[9][23] ), .C(\regs[10][23] ), .D(
        \regs[11][23] ), .S0(n1824), .S1(n1801), .Y(n1695) );
  MX4X1 U2277 ( .A(\regs[8][24] ), .B(\regs[9][24] ), .C(\regs[10][24] ), .D(
        \regs[11][24] ), .S0(n1825), .S1(n1802), .Y(n1705) );
  MX4X1 U2278 ( .A(\regs[8][25] ), .B(\regs[9][25] ), .C(\regs[10][25] ), .D(
        \regs[11][25] ), .S0(n1825), .S1(n1802), .Y(n1715) );
  MX4X1 U2279 ( .A(\regs[8][26] ), .B(\regs[9][26] ), .C(\regs[10][26] ), .D(
        \regs[11][26] ), .S0(n1826), .S1(n1803), .Y(n1725) );
  MX4X1 U2280 ( .A(\regs[8][27] ), .B(\regs[9][27] ), .C(\regs[10][27] ), .D(
        \regs[11][27] ), .S0(n1827), .S1(n1804), .Y(n1735) );
  MX4X1 U2281 ( .A(\regs[8][28] ), .B(\regs[9][28] ), .C(\regs[10][28] ), .D(
        \regs[11][28] ), .S0(n1827), .S1(n1804), .Y(n1745) );
  MX4X1 U2282 ( .A(\regs[8][29] ), .B(\regs[9][29] ), .C(\regs[10][29] ), .D(
        \regs[11][29] ), .S0(n1828), .S1(n1805), .Y(n1755) );
  MX4X1 U2283 ( .A(\regs[8][30] ), .B(\regs[9][30] ), .C(\regs[10][30] ), .D(
        \regs[11][30] ), .S0(n1829), .S1(n1806), .Y(n1765) );
  MX4X1 U2284 ( .A(\regs[8][31] ), .B(\regs[9][31] ), .C(\regs[10][31] ), .D(
        \regs[11][31] ), .S0(n1829), .S1(n1806), .Y(n1775) );
  MX4X1 U2285 ( .A(n1472), .B(n1470), .C(n1471), .D(n1469), .S0(N20), .S1(
        n1783), .Y(n1473) );
  MX4X1 U2286 ( .A(\regs[16][1] ), .B(\regs[17][1] ), .C(\regs[18][1] ), .D(
        \regs[19][1] ), .S0(n1809), .S1(n1786), .Y(n1472) );
  MX4X1 U2287 ( .A(\regs[24][1] ), .B(\regs[25][1] ), .C(\regs[26][1] ), .D(
        \regs[27][1] ), .S0(n1809), .S1(n1786), .Y(n1470) );
  MX4X1 U2288 ( .A(\regs[20][1] ), .B(\regs[21][1] ), .C(\regs[22][1] ), .D(
        \regs[23][1] ), .S0(n1809), .S1(n1786), .Y(n1471) );
  MX4X1 U2289 ( .A(n1482), .B(n1480), .C(n1481), .D(n1479), .S0(n1781), .S1(
        n1783), .Y(n1483) );
  MX4X1 U2290 ( .A(\regs[16][2] ), .B(\regs[17][2] ), .C(\regs[18][2] ), .D(
        \regs[19][2] ), .S0(n1810), .S1(n1787), .Y(n1482) );
  MX4X1 U2291 ( .A(\regs[24][2] ), .B(\regs[25][2] ), .C(\regs[26][2] ), .D(
        \regs[27][2] ), .S0(n1810), .S1(n1787), .Y(n1480) );
  MX4X1 U2292 ( .A(\regs[20][2] ), .B(\regs[21][2] ), .C(\regs[22][2] ), .D(
        \regs[23][2] ), .S0(n1810), .S1(n1787), .Y(n1481) );
  MX4X1 U2293 ( .A(n1492), .B(n1490), .C(n1491), .D(n1489), .S0(n1781), .S1(
        n1783), .Y(n1493) );
  MX4X1 U2294 ( .A(\regs[16][3] ), .B(\regs[17][3] ), .C(\regs[18][3] ), .D(
        \regs[19][3] ), .S0(n1810), .S1(n1787), .Y(n1492) );
  MX4X1 U2295 ( .A(\regs[24][3] ), .B(\regs[25][3] ), .C(\regs[26][3] ), .D(
        \regs[27][3] ), .S0(n1810), .S1(n1787), .Y(n1490) );
  MX4X1 U2296 ( .A(\regs[20][3] ), .B(\regs[21][3] ), .C(\regs[22][3] ), .D(
        \regs[23][3] ), .S0(n1810), .S1(n1787), .Y(n1491) );
  MX4X1 U2297 ( .A(n1502), .B(n1500), .C(n1501), .D(n1499), .S0(n1780), .S1(
        n1783), .Y(n1503) );
  MX4X1 U2298 ( .A(\regs[16][4] ), .B(\regs[17][4] ), .C(\regs[18][4] ), .D(
        \regs[19][4] ), .S0(n1811), .S1(n1788), .Y(n1502) );
  MX4X1 U2299 ( .A(\regs[24][4] ), .B(\regs[25][4] ), .C(\regs[26][4] ), .D(
        \regs[27][4] ), .S0(n1811), .S1(n1788), .Y(n1500) );
  MX4X1 U2300 ( .A(\regs[20][4] ), .B(\regs[21][4] ), .C(\regs[22][4] ), .D(
        \regs[23][4] ), .S0(n1811), .S1(n1788), .Y(n1501) );
  MX4X1 U2301 ( .A(n1512), .B(n1510), .C(n1511), .D(n1509), .S0(n1781), .S1(
        n1783), .Y(n1513) );
  MX4X1 U2302 ( .A(\regs[16][5] ), .B(\regs[17][5] ), .C(\regs[18][5] ), .D(
        \regs[19][5] ), .S0(n1812), .S1(n1789), .Y(n1512) );
  MX4X1 U2303 ( .A(\regs[24][5] ), .B(\regs[25][5] ), .C(\regs[26][5] ), .D(
        \regs[27][5] ), .S0(n1812), .S1(n1789), .Y(n1510) );
  MX4X1 U2304 ( .A(\regs[20][5] ), .B(\regs[21][5] ), .C(\regs[22][5] ), .D(
        \regs[23][5] ), .S0(n1812), .S1(n1789), .Y(n1511) );
  MX4X1 U2305 ( .A(n1522), .B(n1520), .C(n1521), .D(n1519), .S0(n1780), .S1(
        n1783), .Y(n1523) );
  MX4X1 U2306 ( .A(\regs[16][6] ), .B(\regs[17][6] ), .C(\regs[18][6] ), .D(
        \regs[19][6] ), .S0(n1812), .S1(n1789), .Y(n1522) );
  MX4X1 U2307 ( .A(\regs[24][6] ), .B(\regs[25][6] ), .C(\regs[26][6] ), .D(
        \regs[27][6] ), .S0(n1812), .S1(n1789), .Y(n1520) );
  MX4X1 U2308 ( .A(\regs[20][6] ), .B(\regs[21][6] ), .C(\regs[22][6] ), .D(
        \regs[23][6] ), .S0(n1812), .S1(n1789), .Y(n1521) );
  MX4X1 U2309 ( .A(n1532), .B(n1530), .C(n1531), .D(n1529), .S0(n1781), .S1(
        n1783), .Y(n1533) );
  MX4X1 U2310 ( .A(\regs[16][7] ), .B(\regs[17][7] ), .C(\regs[18][7] ), .D(
        \regs[19][7] ), .S0(n1813), .S1(n1790), .Y(n1532) );
  MX4X1 U2311 ( .A(\regs[24][7] ), .B(\regs[25][7] ), .C(\regs[26][7] ), .D(
        \regs[27][7] ), .S0(n1813), .S1(n1790), .Y(n1530) );
  MX4X1 U2312 ( .A(\regs[20][7] ), .B(\regs[21][7] ), .C(\regs[22][7] ), .D(
        \regs[23][7] ), .S0(n1813), .S1(n1790), .Y(n1531) );
  MX4X1 U2313 ( .A(n1542), .B(n1540), .C(n1541), .D(n1539), .S0(n1780), .S1(
        n1783), .Y(n1543) );
  MX4X1 U2314 ( .A(\regs[16][8] ), .B(\regs[17][8] ), .C(\regs[18][8] ), .D(
        \regs[19][8] ), .S0(n1814), .S1(n1791), .Y(n1542) );
  MX4X1 U2315 ( .A(\regs[24][8] ), .B(\regs[25][8] ), .C(\regs[26][8] ), .D(
        \regs[27][8] ), .S0(n1814), .S1(n1791), .Y(n1540) );
  MX4X1 U2316 ( .A(\regs[20][8] ), .B(\regs[21][8] ), .C(\regs[22][8] ), .D(
        \regs[23][8] ), .S0(n1814), .S1(n1791), .Y(n1541) );
  MX4X1 U2317 ( .A(n1552), .B(n1550), .C(n1551), .D(n1549), .S0(N20), .S1(N19), 
        .Y(n1553) );
  MX4X1 U2318 ( .A(\regs[16][9] ), .B(\regs[17][9] ), .C(\regs[18][9] ), .D(
        \regs[19][9] ), .S0(n1814), .S1(n1791), .Y(n1552) );
  MX4X1 U2319 ( .A(\regs[24][9] ), .B(\regs[25][9] ), .C(\regs[26][9] ), .D(
        \regs[27][9] ), .S0(n1814), .S1(n1791), .Y(n1550) );
  MX4X1 U2320 ( .A(\regs[20][9] ), .B(\regs[21][9] ), .C(\regs[22][9] ), .D(
        \regs[23][9] ), .S0(n1814), .S1(n1791), .Y(n1551) );
  MX4X1 U2321 ( .A(n1562), .B(n1560), .C(n1561), .D(n1559), .S0(N20), .S1(N19), 
        .Y(n1563) );
  MX4X1 U2322 ( .A(\regs[16][10] ), .B(\regs[17][10] ), .C(\regs[18][10] ), 
        .D(\regs[19][10] ), .S0(n1815), .S1(n1792), .Y(n1562) );
  MX4X1 U2323 ( .A(\regs[24][10] ), .B(\regs[25][10] ), .C(\regs[26][10] ), 
        .D(\regs[27][10] ), .S0(n1815), .S1(n1792), .Y(n1560) );
  MX4X1 U2324 ( .A(\regs[20][10] ), .B(\regs[21][10] ), .C(\regs[22][10] ), 
        .D(\regs[23][10] ), .S0(n1815), .S1(n1792), .Y(n1561) );
  MX4X1 U2325 ( .A(n1572), .B(n1570), .C(n1571), .D(n1569), .S0(n1781), .S1(
        N19), .Y(n1573) );
  MX4X1 U2326 ( .A(\regs[16][11] ), .B(\regs[17][11] ), .C(\regs[18][11] ), 
        .D(\regs[19][11] ), .S0(n1816), .S1(n1793), .Y(n1572) );
  MX4X1 U2327 ( .A(\regs[24][11] ), .B(\regs[25][11] ), .C(\regs[26][11] ), 
        .D(\regs[27][11] ), .S0(n1816), .S1(n1793), .Y(n1570) );
  MX4X1 U2328 ( .A(\regs[20][11] ), .B(\regs[21][11] ), .C(\regs[22][11] ), 
        .D(\regs[23][11] ), .S0(n1816), .S1(n1793), .Y(n1571) );
  MX4X1 U2329 ( .A(n1582), .B(n1580), .C(n1581), .D(n1579), .S0(N20), .S1(N19), 
        .Y(n1583) );
  MX4X1 U2330 ( .A(\regs[16][12] ), .B(\regs[17][12] ), .C(\regs[18][12] ), 
        .D(\regs[19][12] ), .S0(n1816), .S1(n1793), .Y(n1582) );
  MX4X1 U2331 ( .A(\regs[24][12] ), .B(\regs[25][12] ), .C(\regs[26][12] ), 
        .D(\regs[27][12] ), .S0(n1816), .S1(n1793), .Y(n1580) );
  MX4X1 U2332 ( .A(\regs[20][12] ), .B(\regs[21][12] ), .C(\regs[22][12] ), 
        .D(\regs[23][12] ), .S0(n1816), .S1(n1793), .Y(n1581) );
  MX4X1 U2333 ( .A(n1592), .B(n1590), .C(n1591), .D(n1589), .S0(n1780), .S1(
        N19), .Y(n1593) );
  MX4X1 U2334 ( .A(\regs[16][13] ), .B(\regs[17][13] ), .C(\regs[18][13] ), 
        .D(\regs[19][13] ), .S0(n1817), .S1(n1794), .Y(n1592) );
  MX4X1 U2335 ( .A(\regs[24][13] ), .B(\regs[25][13] ), .C(\regs[26][13] ), 
        .D(\regs[27][13] ), .S0(n1817), .S1(n1794), .Y(n1590) );
  MX4X1 U2336 ( .A(\regs[20][13] ), .B(\regs[21][13] ), .C(\regs[22][13] ), 
        .D(\regs[23][13] ), .S0(n1817), .S1(n1794), .Y(n1591) );
  MX4X1 U2337 ( .A(n1602), .B(n1600), .C(n1601), .D(n1599), .S0(n1780), .S1(
        N19), .Y(n1603) );
  MX4X1 U2338 ( .A(\regs[16][14] ), .B(\regs[17][14] ), .C(\regs[18][14] ), 
        .D(\regs[19][14] ), .S0(n1818), .S1(n1795), .Y(n1602) );
  MX4X1 U2339 ( .A(\regs[24][14] ), .B(\regs[25][14] ), .C(\regs[26][14] ), 
        .D(\regs[27][14] ), .S0(n1818), .S1(n1795), .Y(n1600) );
  MX4X1 U2340 ( .A(\regs[20][14] ), .B(\regs[21][14] ), .C(\regs[22][14] ), 
        .D(\regs[23][14] ), .S0(n1818), .S1(n1795), .Y(n1601) );
  MX4X1 U2341 ( .A(n1612), .B(n1610), .C(n1611), .D(n1609), .S0(n1780), .S1(
        N19), .Y(n1613) );
  MX4X1 U2342 ( .A(\regs[16][15] ), .B(\regs[17][15] ), .C(\regs[18][15] ), 
        .D(\regs[19][15] ), .S0(n1818), .S1(n1795), .Y(n1612) );
  MX4X1 U2343 ( .A(\regs[24][15] ), .B(\regs[25][15] ), .C(\regs[26][15] ), 
        .D(\regs[27][15] ), .S0(n1818), .S1(n1795), .Y(n1610) );
  MX4X1 U2344 ( .A(\regs[20][15] ), .B(\regs[21][15] ), .C(\regs[22][15] ), 
        .D(\regs[23][15] ), .S0(n1818), .S1(n1795), .Y(n1611) );
  MX4X1 U2345 ( .A(n1622), .B(n1620), .C(n1621), .D(n1619), .S0(n1780), .S1(
        N19), .Y(n1623) );
  MX4X1 U2346 ( .A(\regs[16][16] ), .B(\regs[17][16] ), .C(\regs[18][16] ), 
        .D(\regs[19][16] ), .S0(n1819), .S1(n1796), .Y(n1622) );
  MX4X1 U2347 ( .A(\regs[24][16] ), .B(\regs[25][16] ), .C(\regs[26][16] ), 
        .D(\regs[27][16] ), .S0(n1819), .S1(n1796), .Y(n1620) );
  MX4X1 U2348 ( .A(\regs[20][16] ), .B(\regs[21][16] ), .C(\regs[22][16] ), 
        .D(\regs[23][16] ), .S0(n1819), .S1(n1796), .Y(n1621) );
  MX4X1 U2349 ( .A(n1632), .B(n1630), .C(n1631), .D(n1629), .S0(n1780), .S1(
        n1783), .Y(n1633) );
  MX4X1 U2350 ( .A(\regs[16][17] ), .B(\regs[17][17] ), .C(\regs[18][17] ), 
        .D(\regs[19][17] ), .S0(n1820), .S1(n1797), .Y(n1632) );
  MX4X1 U2351 ( .A(\regs[24][17] ), .B(\regs[25][17] ), .C(\regs[26][17] ), 
        .D(\regs[27][17] ), .S0(n1820), .S1(n1797), .Y(n1630) );
  MX4X1 U2352 ( .A(\regs[20][17] ), .B(\regs[21][17] ), .C(\regs[22][17] ), 
        .D(\regs[23][17] ), .S0(n1820), .S1(n1797), .Y(n1631) );
  MX4X1 U2353 ( .A(n1642), .B(n1640), .C(n1641), .D(n1639), .S0(n1780), .S1(
        N19), .Y(n1643) );
  MX4X1 U2354 ( .A(\regs[16][18] ), .B(\regs[17][18] ), .C(\regs[18][18] ), 
        .D(\regs[19][18] ), .S0(n1820), .S1(n1797), .Y(n1642) );
  MX4X1 U2355 ( .A(\regs[24][18] ), .B(\regs[25][18] ), .C(\regs[26][18] ), 
        .D(\regs[27][18] ), .S0(n1820), .S1(n1797), .Y(n1640) );
  MX4X1 U2356 ( .A(\regs[20][18] ), .B(\regs[21][18] ), .C(\regs[22][18] ), 
        .D(\regs[23][18] ), .S0(n1820), .S1(n1797), .Y(n1641) );
  MX4X1 U2357 ( .A(n1652), .B(n1650), .C(n1651), .D(n1649), .S0(n1780), .S1(
        N19), .Y(n1653) );
  MX4X1 U2358 ( .A(\regs[16][19] ), .B(\regs[17][19] ), .C(\regs[18][19] ), 
        .D(\regs[19][19] ), .S0(n1821), .S1(n1798), .Y(n1652) );
  MX4X1 U2359 ( .A(\regs[24][19] ), .B(\regs[25][19] ), .C(\regs[26][19] ), 
        .D(\regs[27][19] ), .S0(n1821), .S1(n1798), .Y(n1650) );
  MX4X1 U2360 ( .A(\regs[20][19] ), .B(\regs[21][19] ), .C(\regs[22][19] ), 
        .D(\regs[23][19] ), .S0(n1821), .S1(n1798), .Y(n1651) );
  MX4X1 U2361 ( .A(n1662), .B(n1660), .C(n1661), .D(n1659), .S0(n1781), .S1(
        N19), .Y(n1663) );
  MX4X1 U2362 ( .A(\regs[16][20] ), .B(\regs[17][20] ), .C(\regs[18][20] ), 
        .D(\regs[19][20] ), .S0(n1822), .S1(n1799), .Y(n1662) );
  MX4X1 U2363 ( .A(\regs[24][20] ), .B(\regs[25][20] ), .C(\regs[26][20] ), 
        .D(\regs[27][20] ), .S0(n1822), .S1(n1799), .Y(n1660) );
  MX4X1 U2364 ( .A(\regs[20][20] ), .B(\regs[21][20] ), .C(\regs[22][20] ), 
        .D(\regs[23][20] ), .S0(n1822), .S1(n1799), .Y(n1661) );
  MX4X1 U2365 ( .A(n1672), .B(n1670), .C(n1671), .D(n1669), .S0(n1781), .S1(
        N19), .Y(n1673) );
  MX4X1 U2366 ( .A(\regs[16][21] ), .B(\regs[17][21] ), .C(\regs[18][21] ), 
        .D(\regs[19][21] ), .S0(n1822), .S1(n1799), .Y(n1672) );
  MX4X1 U2367 ( .A(\regs[24][21] ), .B(\regs[25][21] ), .C(\regs[26][21] ), 
        .D(\regs[27][21] ), .S0(n1822), .S1(n1799), .Y(n1670) );
  MX4X1 U2368 ( .A(\regs[20][21] ), .B(\regs[21][21] ), .C(\regs[22][21] ), 
        .D(\regs[23][21] ), .S0(n1822), .S1(n1799), .Y(n1671) );
  MX4X1 U2369 ( .A(n1682), .B(n1680), .C(n1681), .D(n1679), .S0(n1781), .S1(
        N19), .Y(n1683) );
  MX4X1 U2370 ( .A(\regs[16][22] ), .B(\regs[17][22] ), .C(\regs[18][22] ), 
        .D(\regs[19][22] ), .S0(n1823), .S1(n1800), .Y(n1682) );
  MX4X1 U2371 ( .A(\regs[24][22] ), .B(\regs[25][22] ), .C(\regs[26][22] ), 
        .D(\regs[27][22] ), .S0(n1823), .S1(n1800), .Y(n1680) );
  MX4X1 U2372 ( .A(\regs[20][22] ), .B(\regs[21][22] ), .C(\regs[22][22] ), 
        .D(\regs[23][22] ), .S0(n1823), .S1(n1800), .Y(n1681) );
  MX4X1 U2373 ( .A(n1692), .B(n1690), .C(n1691), .D(n1689), .S0(n1781), .S1(
        N19), .Y(n1693) );
  MX4X1 U2374 ( .A(\regs[16][23] ), .B(\regs[17][23] ), .C(\regs[18][23] ), 
        .D(\regs[19][23] ), .S0(n1824), .S1(n1801), .Y(n1692) );
  MX4X1 U2375 ( .A(\regs[24][23] ), .B(\regs[25][23] ), .C(\regs[26][23] ), 
        .D(\regs[27][23] ), .S0(n1824), .S1(n1801), .Y(n1690) );
  MX4X1 U2376 ( .A(\regs[20][23] ), .B(\regs[21][23] ), .C(\regs[22][23] ), 
        .D(\regs[23][23] ), .S0(n1824), .S1(n1801), .Y(n1691) );
  MX4X1 U2377 ( .A(n1702), .B(n1700), .C(n1701), .D(n1699), .S0(n1781), .S1(
        n1783), .Y(n1703) );
  MX4X1 U2378 ( .A(\regs[16][24] ), .B(\regs[17][24] ), .C(\regs[18][24] ), 
        .D(\regs[19][24] ), .S0(n1824), .S1(n1801), .Y(n1702) );
  MX4X1 U2379 ( .A(\regs[24][24] ), .B(\regs[25][24] ), .C(\regs[26][24] ), 
        .D(\regs[27][24] ), .S0(n1824), .S1(n1801), .Y(n1700) );
  MX4X1 U2380 ( .A(\regs[20][24] ), .B(\regs[21][24] ), .C(\regs[22][24] ), 
        .D(\regs[23][24] ), .S0(n1824), .S1(n1801), .Y(n1701) );
  MX4X1 U2381 ( .A(n1712), .B(n1710), .C(n1711), .D(n1709), .S0(n1781), .S1(
        N19), .Y(n1713) );
  MX4X1 U2382 ( .A(\regs[16][25] ), .B(\regs[17][25] ), .C(\regs[18][25] ), 
        .D(\regs[19][25] ), .S0(n1825), .S1(n1802), .Y(n1712) );
  MX4X1 U2383 ( .A(\regs[24][25] ), .B(\regs[25][25] ), .C(\regs[26][25] ), 
        .D(\regs[27][25] ), .S0(n1825), .S1(n1802), .Y(n1710) );
  MX4X1 U2384 ( .A(\regs[20][25] ), .B(\regs[21][25] ), .C(\regs[22][25] ), 
        .D(\regs[23][25] ), .S0(n1825), .S1(n1802), .Y(n1711) );
  MX4X1 U2385 ( .A(n1722), .B(n1720), .C(n1721), .D(n1719), .S0(n1781), .S1(
        N19), .Y(n1723) );
  MX4X1 U2386 ( .A(\regs[16][26] ), .B(\regs[17][26] ), .C(\regs[18][26] ), 
        .D(\regs[19][26] ), .S0(n1826), .S1(n1803), .Y(n1722) );
  MX4X1 U2387 ( .A(\regs[24][26] ), .B(\regs[25][26] ), .C(\regs[26][26] ), 
        .D(\regs[27][26] ), .S0(n1826), .S1(n1803), .Y(n1720) );
  MX4X1 U2388 ( .A(\regs[20][26] ), .B(\regs[21][26] ), .C(\regs[22][26] ), 
        .D(\regs[23][26] ), .S0(n1826), .S1(n1803), .Y(n1721) );
  MX4X1 U2389 ( .A(n1732), .B(n1730), .C(n1731), .D(n1729), .S0(n1780), .S1(
        N19), .Y(n1733) );
  MX4X1 U2390 ( .A(\regs[16][27] ), .B(\regs[17][27] ), .C(\regs[18][27] ), 
        .D(\regs[19][27] ), .S0(n1826), .S1(n1803), .Y(n1732) );
  MX4X1 U2391 ( .A(\regs[24][27] ), .B(\regs[25][27] ), .C(\regs[26][27] ), 
        .D(\regs[27][27] ), .S0(n1826), .S1(n1803), .Y(n1730) );
  MX4X1 U2392 ( .A(\regs[20][27] ), .B(\regs[21][27] ), .C(\regs[22][27] ), 
        .D(\regs[23][27] ), .S0(n1826), .S1(n1803), .Y(n1731) );
  MX4X1 U2393 ( .A(n1742), .B(n1740), .C(n1741), .D(n1739), .S0(n1780), .S1(
        N19), .Y(n1743) );
  MX4X1 U2394 ( .A(\regs[16][28] ), .B(\regs[17][28] ), .C(\regs[18][28] ), 
        .D(\regs[19][28] ), .S0(n1827), .S1(n1804), .Y(n1742) );
  MX4X1 U2395 ( .A(\regs[24][28] ), .B(\regs[25][28] ), .C(\regs[26][28] ), 
        .D(\regs[27][28] ), .S0(n1827), .S1(n1804), .Y(n1740) );
  MX4X1 U2396 ( .A(\regs[20][28] ), .B(\regs[21][28] ), .C(\regs[22][28] ), 
        .D(\regs[23][28] ), .S0(n1827), .S1(n1804), .Y(n1741) );
  MX4X1 U2397 ( .A(n1752), .B(n1750), .C(n1751), .D(n1749), .S0(N20), .S1(N19), 
        .Y(n1753) );
  MX4X1 U2398 ( .A(\regs[16][29] ), .B(\regs[17][29] ), .C(\regs[18][29] ), 
        .D(\regs[19][29] ), .S0(n1828), .S1(n1805), .Y(n1752) );
  MX4X1 U2399 ( .A(\regs[24][29] ), .B(\regs[25][29] ), .C(\regs[26][29] ), 
        .D(\regs[27][29] ), .S0(n1828), .S1(n1805), .Y(n1750) );
  MX4X1 U2400 ( .A(\regs[20][29] ), .B(\regs[21][29] ), .C(\regs[22][29] ), 
        .D(\regs[23][29] ), .S0(n1828), .S1(n1805), .Y(n1751) );
  MX4X1 U2401 ( .A(n1762), .B(n1760), .C(n1761), .D(n1759), .S0(N20), .S1(
        n1783), .Y(n1763) );
  MX4X1 U2402 ( .A(\regs[16][30] ), .B(\regs[17][30] ), .C(\regs[18][30] ), 
        .D(\regs[19][30] ), .S0(n1828), .S1(n1805), .Y(n1762) );
  MX4X1 U2403 ( .A(\regs[24][30] ), .B(\regs[25][30] ), .C(\regs[26][30] ), 
        .D(\regs[27][30] ), .S0(n1828), .S1(n1805), .Y(n1760) );
  MX4X1 U2404 ( .A(\regs[20][30] ), .B(\regs[21][30] ), .C(\regs[22][30] ), 
        .D(\regs[23][30] ), .S0(n1828), .S1(n1805), .Y(n1761) );
  MX4X1 U2405 ( .A(n1772), .B(n1770), .C(n1771), .D(n1769), .S0(N20), .S1(
        n1783), .Y(n1773) );
  MX4X1 U2406 ( .A(\regs[16][31] ), .B(\regs[17][31] ), .C(\regs[18][31] ), 
        .D(\regs[19][31] ), .S0(n1829), .S1(n1806), .Y(n1772) );
  MX4X1 U2407 ( .A(\regs[24][31] ), .B(\regs[25][31] ), .C(\regs[26][31] ), 
        .D(\regs[27][31] ), .S0(n1829), .S1(n1806), .Y(n1770) );
  MX4X1 U2408 ( .A(\regs[20][31] ), .B(\regs[21][31] ), .C(\regs[22][31] ), 
        .D(\regs[23][31] ), .S0(n1829), .S1(n1806), .Y(n1771) );
  NOR2X1 U2409 ( .A(write_addr[0]), .B(write_addr[1]), .Y(n35) );
  NOR2X1 U2410 ( .A(n83), .B(write_addr[1]), .Y(n38) );
  AND2X2 U2411 ( .A(write_addr[1]), .B(n83), .Y(n40) );
  AND2X2 U2412 ( .A(write_addr[1]), .B(write_addr[0]), .Y(n42) );
  NOR2BX1 U2413 ( .AN(reg_rw), .B(write_addr[4]), .Y(n43) );
  NOR2X1 U2414 ( .A(write_addr[2]), .B(write_addr[3]), .Y(n44) );
  NOR2X1 U2415 ( .A(n74), .B(write_addr[3]), .Y(n50) );
  INVX1 U2416 ( .A(write_addr[0]), .Y(n83) );
  INVX1 U2417 ( .A(write_addr[2]), .Y(n74) );
  AND2X2 U2418 ( .A(write_addr[4]), .B(reg_rw), .Y(n68) );
  AND2X2 U2419 ( .A(write_addr[3]), .B(n74), .Y(n56) );
  AND2X2 U2420 ( .A(write_addr[3]), .B(write_addr[2]), .Y(n62) );
endmodule


module IFID ( pc_out, inst_out, pc_in, inst_in, clk, rst, flush, stall );
  output [31:0] pc_out;
  output [31:0] inst_out;
  input [31:0] pc_in;
  input [31:0] inst_in;
  input clk, rst, flush, stall;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n1, n132, n133,
         n134;

  DFFRHQX1 \inst_out_reg[31]  ( .D(n99), .CK(clk), .RN(rst), .Q(inst_out[31])
         );
  DFFRHQX1 \pc_out_reg[31]  ( .D(n131), .CK(clk), .RN(rst), .Q(pc_out[31]) );
  DFFRHQX1 \pc_out_reg[30]  ( .D(n130), .CK(clk), .RN(rst), .Q(pc_out[30]) );
  DFFRHQX1 \pc_out_reg[29]  ( .D(n129), .CK(clk), .RN(rst), .Q(pc_out[29]) );
  DFFRHQX1 \pc_out_reg[28]  ( .D(n128), .CK(clk), .RN(rst), .Q(pc_out[28]) );
  DFFRHQX1 \pc_out_reg[27]  ( .D(n127), .CK(clk), .RN(rst), .Q(pc_out[27]) );
  DFFRHQX1 \pc_out_reg[26]  ( .D(n126), .CK(clk), .RN(rst), .Q(pc_out[26]) );
  DFFRHQX1 \pc_out_reg[25]  ( .D(n125), .CK(clk), .RN(rst), .Q(pc_out[25]) );
  DFFRHQX1 \pc_out_reg[24]  ( .D(n124), .CK(clk), .RN(rst), .Q(pc_out[24]) );
  DFFRHQX1 \pc_out_reg[23]  ( .D(n123), .CK(clk), .RN(rst), .Q(pc_out[23]) );
  DFFRHQX1 \pc_out_reg[22]  ( .D(n122), .CK(clk), .RN(rst), .Q(pc_out[22]) );
  DFFRHQX1 \pc_out_reg[21]  ( .D(n121), .CK(clk), .RN(rst), .Q(pc_out[21]) );
  DFFRHQX1 \pc_out_reg[20]  ( .D(n120), .CK(clk), .RN(rst), .Q(pc_out[20]) );
  DFFRHQX1 \pc_out_reg[19]  ( .D(n119), .CK(clk), .RN(rst), .Q(pc_out[19]) );
  DFFRHQX1 \pc_out_reg[18]  ( .D(n118), .CK(clk), .RN(rst), .Q(pc_out[18]) );
  DFFRHQX1 \pc_out_reg[17]  ( .D(n117), .CK(clk), .RN(rst), .Q(pc_out[17]) );
  DFFRHQX1 \pc_out_reg[16]  ( .D(n116), .CK(clk), .RN(rst), .Q(pc_out[16]) );
  DFFRHQX1 \pc_out_reg[15]  ( .D(n115), .CK(clk), .RN(rst), .Q(pc_out[15]) );
  DFFRHQX1 \inst_out_reg[24]  ( .D(n92), .CK(clk), .RN(rst), .Q(inst_out[24])
         );
  DFFRHQX1 \inst_out_reg[23]  ( .D(n91), .CK(clk), .RN(rst), .Q(inst_out[23])
         );
  DFFRHQX1 \inst_out_reg[22]  ( .D(n90), .CK(clk), .RN(rst), .Q(inst_out[22])
         );
  DFFRHQX1 \inst_out_reg[21]  ( .D(n89), .CK(clk), .RN(rst), .Q(inst_out[21])
         );
  DFFRHQX1 \inst_out_reg[20]  ( .D(n88), .CK(clk), .RN(rst), .Q(inst_out[20])
         );
  DFFRHQX1 \inst_out_reg[19]  ( .D(n87), .CK(clk), .RN(rst), .Q(inst_out[19])
         );
  DFFRHQX1 \inst_out_reg[18]  ( .D(n86), .CK(clk), .RN(rst), .Q(inst_out[18])
         );
  DFFRHQX1 \inst_out_reg[17]  ( .D(n85), .CK(clk), .RN(rst), .Q(inst_out[17])
         );
  DFFRHQX1 \inst_out_reg[16]  ( .D(n84), .CK(clk), .RN(rst), .Q(inst_out[16])
         );
  DFFRHQX1 \inst_out_reg[15]  ( .D(n83), .CK(clk), .RN(rst), .Q(inst_out[15])
         );
  DFFRHQX1 \pc_out_reg[14]  ( .D(n114), .CK(clk), .RN(rst), .Q(pc_out[14]) );
  DFFRHQX1 \pc_out_reg[13]  ( .D(n113), .CK(clk), .RN(rst), .Q(pc_out[13]) );
  DFFRHQX1 \pc_out_reg[12]  ( .D(n112), .CK(clk), .RN(rst), .Q(pc_out[12]) );
  DFFRHQX1 \pc_out_reg[11]  ( .D(n111), .CK(clk), .RN(rst), .Q(pc_out[11]) );
  DFFRHQX1 \pc_out_reg[10]  ( .D(n110), .CK(clk), .RN(rst), .Q(pc_out[10]) );
  DFFRHQX1 \pc_out_reg[9]  ( .D(n109), .CK(clk), .RN(rst), .Q(pc_out[9]) );
  DFFRHQX1 \pc_out_reg[8]  ( .D(n108), .CK(clk), .RN(rst), .Q(pc_out[8]) );
  DFFRHQX1 \pc_out_reg[7]  ( .D(n107), .CK(clk), .RN(rst), .Q(pc_out[7]) );
  DFFRHQX1 \pc_out_reg[6]  ( .D(n106), .CK(clk), .RN(rst), .Q(pc_out[6]) );
  DFFRHQX1 \pc_out_reg[5]  ( .D(n105), .CK(clk), .RN(rst), .Q(pc_out[5]) );
  DFFRHQX1 \inst_out_reg[9]  ( .D(n77), .CK(clk), .RN(rst), .Q(inst_out[9]) );
  DFFRHQX1 \inst_out_reg[8]  ( .D(n76), .CK(clk), .RN(rst), .Q(inst_out[8]) );
  DFFRHQX1 \inst_out_reg[7]  ( .D(n75), .CK(clk), .RN(rst), .Q(inst_out[7]) );
  DFFRHQX1 \inst_out_reg[6]  ( .D(n74), .CK(clk), .RN(rst), .Q(inst_out[6]) );
  DFFRHQX1 \inst_out_reg[5]  ( .D(n73), .CK(clk), .RN(rst), .Q(inst_out[5]) );
  DFFRHQX1 \pc_out_reg[0]  ( .D(n100), .CK(clk), .RN(rst), .Q(pc_out[0]) );
  DFFRHQX1 \inst_out_reg[14]  ( .D(n82), .CK(clk), .RN(rst), .Q(inst_out[14])
         );
  DFFRHQX1 \inst_out_reg[13]  ( .D(n81), .CK(clk), .RN(rst), .Q(inst_out[13])
         );
  DFFRHQX1 \inst_out_reg[12]  ( .D(n80), .CK(clk), .RN(rst), .Q(inst_out[12])
         );
  DFFRHQX1 \inst_out_reg[11]  ( .D(n79), .CK(clk), .RN(rst), .Q(inst_out[11])
         );
  DFFRHQX1 \inst_out_reg[10]  ( .D(n78), .CK(clk), .RN(rst), .Q(inst_out[10])
         );
  DFFRHQX1 \pc_out_reg[4]  ( .D(n104), .CK(clk), .RN(rst), .Q(pc_out[4]) );
  DFFRHQX1 \pc_out_reg[3]  ( .D(n103), .CK(clk), .RN(rst), .Q(pc_out[3]) );
  DFFRHQX1 \pc_out_reg[2]  ( .D(n102), .CK(clk), .RN(rst), .Q(pc_out[2]) );
  DFFRHQX1 \pc_out_reg[1]  ( .D(n101), .CK(clk), .RN(rst), .Q(pc_out[1]) );
  DFFRHQX1 \inst_out_reg[4]  ( .D(n72), .CK(clk), .RN(rst), .Q(inst_out[4]) );
  DFFRHQX1 \inst_out_reg[2]  ( .D(n70), .CK(clk), .RN(rst), .Q(inst_out[2]) );
  DFFRHQX1 \inst_out_reg[3]  ( .D(n71), .CK(clk), .RN(rst), .Q(inst_out[3]) );
  DFFRHQX1 \inst_out_reg[0]  ( .D(n68), .CK(clk), .RN(rst), .Q(inst_out[0]) );
  DFFRHQX1 \inst_out_reg[1]  ( .D(n69), .CK(clk), .RN(rst), .Q(inst_out[1]) );
  DFFRHQX1 \inst_out_reg[30]  ( .D(n98), .CK(clk), .RN(rst), .Q(inst_out[30])
         );
  DFFRHQX1 \inst_out_reg[27]  ( .D(n95), .CK(clk), .RN(rst), .Q(inst_out[27])
         );
  DFFRHQX1 \inst_out_reg[29]  ( .D(n97), .CK(clk), .RN(rst), .Q(inst_out[29])
         );
  DFFRHQX1 \inst_out_reg[25]  ( .D(n93), .CK(clk), .RN(rst), .Q(inst_out[25])
         );
  DFFRHQX1 \inst_out_reg[26]  ( .D(n94), .CK(clk), .RN(rst), .Q(inst_out[26])
         );
  DFFRHQX1 \inst_out_reg[28]  ( .D(n96), .CK(clk), .RN(rst), .Q(inst_out[28])
         );
  INVX1 U2 ( .A(n134), .Y(n133) );
  INVX1 U3 ( .A(n132), .Y(n1) );
  INVX1 U4 ( .A(n3), .Y(n134) );
  NOR2X1 U5 ( .A(n4), .B(flush), .Y(n3) );
  INVX1 U6 ( .A(n4), .Y(n132) );
  NOR2BX1 U7 ( .AN(stall), .B(flush), .Y(n4) );
  INVX1 U8 ( .A(n2), .Y(n68) );
  AOI22X1 U9 ( .A0(inst_in[0]), .A1(n3), .B0(inst_out[0]), .B1(n1), .Y(n2) );
  INVX1 U10 ( .A(n9), .Y(n73) );
  AOI22X1 U11 ( .A0(inst_in[5]), .A1(n3), .B0(inst_out[5]), .B1(n1), .Y(n9) );
  INVX1 U12 ( .A(n10), .Y(n74) );
  AOI22X1 U13 ( .A0(inst_in[6]), .A1(n3), .B0(inst_out[6]), .B1(n1), .Y(n10)
         );
  INVX1 U14 ( .A(n11), .Y(n75) );
  AOI22X1 U15 ( .A0(inst_in[7]), .A1(n3), .B0(inst_out[7]), .B1(n1), .Y(n11)
         );
  INVX1 U16 ( .A(n12), .Y(n76) );
  AOI22X1 U17 ( .A0(inst_in[8]), .A1(n3), .B0(inst_out[8]), .B1(n1), .Y(n12)
         );
  INVX1 U18 ( .A(n13), .Y(n77) );
  AOI22X1 U19 ( .A0(inst_in[9]), .A1(n133), .B0(inst_out[9]), .B1(n1), .Y(n13)
         );
  INVX1 U20 ( .A(n31), .Y(n95) );
  AOI22X1 U21 ( .A0(inst_in[27]), .A1(n3), .B0(inst_out[27]), .B1(n1), .Y(n31)
         );
  INVX1 U22 ( .A(n34), .Y(n98) );
  AOI22X1 U23 ( .A0(inst_in[30]), .A1(n3), .B0(inst_out[30]), .B1(n1), .Y(n34)
         );
  INVX1 U24 ( .A(n35), .Y(n99) );
  AOI22X1 U25 ( .A0(inst_in[31]), .A1(n3), .B0(inst_out[31]), .B1(n1), .Y(n35)
         );
  INVX1 U26 ( .A(n37), .Y(n101) );
  AOI22X1 U27 ( .A0(pc_in[1]), .A1(n3), .B0(pc_out[1]), .B1(n1), .Y(n37) );
  INVX1 U28 ( .A(n38), .Y(n102) );
  AOI22X1 U29 ( .A0(pc_in[2]), .A1(n3), .B0(pc_out[2]), .B1(n1), .Y(n38) );
  INVX1 U30 ( .A(n39), .Y(n103) );
  AOI22X1 U31 ( .A0(pc_in[3]), .A1(n3), .B0(pc_out[3]), .B1(n1), .Y(n39) );
  INVX1 U32 ( .A(n40), .Y(n104) );
  AOI22X1 U33 ( .A0(pc_in[4]), .A1(n133), .B0(pc_out[4]), .B1(n1), .Y(n40) );
  INVX1 U34 ( .A(n41), .Y(n105) );
  AOI22X1 U35 ( .A0(pc_in[5]), .A1(n133), .B0(pc_out[5]), .B1(n1), .Y(n41) );
  INVX1 U36 ( .A(n42), .Y(n106) );
  AOI22X1 U37 ( .A0(pc_in[6]), .A1(n133), .B0(pc_out[6]), .B1(n1), .Y(n42) );
  INVX1 U38 ( .A(n43), .Y(n107) );
  AOI22X1 U39 ( .A0(pc_in[7]), .A1(n133), .B0(pc_out[7]), .B1(n1), .Y(n43) );
  INVX1 U40 ( .A(n44), .Y(n108) );
  AOI22X1 U41 ( .A0(pc_in[8]), .A1(n133), .B0(pc_out[8]), .B1(n1), .Y(n44) );
  INVX1 U42 ( .A(n45), .Y(n109) );
  AOI22X1 U43 ( .A0(pc_in[9]), .A1(n133), .B0(pc_out[9]), .B1(n1), .Y(n45) );
  INVX1 U44 ( .A(n46), .Y(n110) );
  AOI22X1 U45 ( .A0(pc_in[10]), .A1(n133), .B0(pc_out[10]), .B1(n1), .Y(n46)
         );
  INVX1 U46 ( .A(n47), .Y(n111) );
  AOI22X1 U47 ( .A0(pc_in[11]), .A1(n133), .B0(pc_out[11]), .B1(n1), .Y(n47)
         );
  INVX1 U48 ( .A(n48), .Y(n112) );
  AOI22X1 U49 ( .A0(pc_in[12]), .A1(n133), .B0(pc_out[12]), .B1(n1), .Y(n48)
         );
  INVX1 U50 ( .A(n49), .Y(n113) );
  AOI22X1 U51 ( .A0(pc_in[13]), .A1(n133), .B0(pc_out[13]), .B1(n1), .Y(n49)
         );
  INVX1 U52 ( .A(n50), .Y(n114) );
  AOI22X1 U53 ( .A0(pc_in[14]), .A1(n133), .B0(pc_out[14]), .B1(n1), .Y(n50)
         );
  INVX1 U54 ( .A(n51), .Y(n115) );
  AOI22X1 U55 ( .A0(pc_in[15]), .A1(n133), .B0(pc_out[15]), .B1(n1), .Y(n51)
         );
  INVX1 U56 ( .A(n52), .Y(n116) );
  AOI22X1 U57 ( .A0(pc_in[16]), .A1(n3), .B0(pc_out[16]), .B1(n1), .Y(n52) );
  INVX1 U58 ( .A(n53), .Y(n117) );
  AOI22X1 U59 ( .A0(pc_in[17]), .A1(n3), .B0(pc_out[17]), .B1(n1), .Y(n53) );
  INVX1 U60 ( .A(n54), .Y(n118) );
  AOI22X1 U61 ( .A0(pc_in[18]), .A1(n3), .B0(pc_out[18]), .B1(n1), .Y(n54) );
  INVX1 U62 ( .A(n55), .Y(n119) );
  AOI22X1 U63 ( .A0(pc_in[19]), .A1(n133), .B0(pc_out[19]), .B1(n1), .Y(n55)
         );
  INVX1 U64 ( .A(n56), .Y(n120) );
  AOI22X1 U65 ( .A0(pc_in[20]), .A1(n3), .B0(pc_out[20]), .B1(n1), .Y(n56) );
  INVX1 U66 ( .A(n57), .Y(n121) );
  AOI22X1 U67 ( .A0(pc_in[21]), .A1(n3), .B0(pc_out[21]), .B1(n1), .Y(n57) );
  INVX1 U68 ( .A(n58), .Y(n122) );
  AOI22X1 U69 ( .A0(pc_in[22]), .A1(n3), .B0(pc_out[22]), .B1(n1), .Y(n58) );
  INVX1 U70 ( .A(n59), .Y(n123) );
  AOI22X1 U71 ( .A0(pc_in[23]), .A1(n133), .B0(pc_out[23]), .B1(n1), .Y(n59)
         );
  INVX1 U72 ( .A(n60), .Y(n124) );
  AOI22X1 U73 ( .A0(pc_in[24]), .A1(n3), .B0(pc_out[24]), .B1(n1), .Y(n60) );
  INVX1 U74 ( .A(n61), .Y(n125) );
  AOI22X1 U75 ( .A0(pc_in[25]), .A1(n133), .B0(pc_out[25]), .B1(n1), .Y(n61)
         );
  INVX1 U76 ( .A(n62), .Y(n126) );
  AOI22X1 U77 ( .A0(pc_in[26]), .A1(n3), .B0(pc_out[26]), .B1(n1), .Y(n62) );
  INVX1 U78 ( .A(n63), .Y(n127) );
  AOI22X1 U79 ( .A0(pc_in[27]), .A1(n3), .B0(pc_out[27]), .B1(n1), .Y(n63) );
  INVX1 U80 ( .A(n64), .Y(n128) );
  AOI22X1 U81 ( .A0(pc_in[28]), .A1(n3), .B0(pc_out[28]), .B1(n1), .Y(n64) );
  INVX1 U82 ( .A(n65), .Y(n129) );
  AOI22X1 U83 ( .A0(pc_in[29]), .A1(n3), .B0(pc_out[29]), .B1(n1), .Y(n65) );
  INVX1 U84 ( .A(n66), .Y(n130) );
  AOI22X1 U85 ( .A0(pc_in[30]), .A1(n3), .B0(pc_out[30]), .B1(n1), .Y(n66) );
  INVX1 U86 ( .A(n67), .Y(n131) );
  AOI22X1 U87 ( .A0(pc_in[31]), .A1(n3), .B0(pc_out[31]), .B1(n1), .Y(n67) );
  INVX1 U88 ( .A(n5), .Y(n69) );
  AOI22X1 U89 ( .A0(inst_in[1]), .A1(n3), .B0(inst_out[1]), .B1(n1), .Y(n5) );
  INVX1 U90 ( .A(n7), .Y(n71) );
  AOI22X1 U91 ( .A0(inst_in[3]), .A1(n3), .B0(inst_out[3]), .B1(n1), .Y(n7) );
  INVX1 U92 ( .A(n32), .Y(n96) );
  AOI22X1 U93 ( .A0(inst_in[28]), .A1(n133), .B0(inst_out[28]), .B1(n1), .Y(
        n32) );
  INVX1 U94 ( .A(n6), .Y(n70) );
  AOI22X1 U95 ( .A0(inst_in[2]), .A1(n3), .B0(inst_out[2]), .B1(n1), .Y(n6) );
  INVX1 U96 ( .A(n30), .Y(n94) );
  AOI22X1 U97 ( .A0(inst_in[26]), .A1(n133), .B0(inst_out[26]), .B1(n1), .Y(
        n30) );
  INVX1 U98 ( .A(n8), .Y(n72) );
  AOI22X1 U99 ( .A0(inst_in[4]), .A1(n133), .B0(inst_out[4]), .B1(n1), .Y(n8)
         );
  INVX1 U100 ( .A(n14), .Y(n78) );
  AOI22X1 U101 ( .A0(inst_in[10]), .A1(n3), .B0(inst_out[10]), .B1(n1), .Y(n14) );
  INVX1 U102 ( .A(n15), .Y(n79) );
  AOI22X1 U103 ( .A0(inst_in[11]), .A1(n3), .B0(inst_out[11]), .B1(n1), .Y(n15) );
  INVX1 U104 ( .A(n16), .Y(n80) );
  AOI22X1 U105 ( .A0(inst_in[12]), .A1(n3), .B0(inst_out[12]), .B1(n1), .Y(n16) );
  INVX1 U106 ( .A(n17), .Y(n81) );
  AOI22X1 U107 ( .A0(inst_in[13]), .A1(n3), .B0(inst_out[13]), .B1(n1), .Y(n17) );
  INVX1 U108 ( .A(n18), .Y(n82) );
  AOI22X1 U109 ( .A0(inst_in[14]), .A1(n3), .B0(inst_out[14]), .B1(n1), .Y(n18) );
  INVX1 U110 ( .A(n19), .Y(n83) );
  AOI22X1 U111 ( .A0(inst_in[15]), .A1(n3), .B0(inst_out[15]), .B1(n1), .Y(n19) );
  INVX1 U112 ( .A(n20), .Y(n84) );
  AOI22X1 U113 ( .A0(inst_in[16]), .A1(n3), .B0(inst_out[16]), .B1(n1), .Y(n20) );
  INVX1 U114 ( .A(n21), .Y(n85) );
  AOI22X1 U115 ( .A0(inst_in[17]), .A1(n133), .B0(inst_out[17]), .B1(n1), .Y(
        n21) );
  INVX1 U116 ( .A(n22), .Y(n86) );
  AOI22X1 U117 ( .A0(inst_in[18]), .A1(n3), .B0(inst_out[18]), .B1(n1), .Y(n22) );
  INVX1 U118 ( .A(n23), .Y(n87) );
  AOI22X1 U119 ( .A0(inst_in[19]), .A1(n3), .B0(inst_out[19]), .B1(n1), .Y(n23) );
  INVX1 U120 ( .A(n24), .Y(n88) );
  AOI22X1 U121 ( .A0(inst_in[20]), .A1(n3), .B0(inst_out[20]), .B1(n1), .Y(n24) );
  INVX1 U122 ( .A(n25), .Y(n89) );
  AOI22X1 U123 ( .A0(inst_in[21]), .A1(n133), .B0(inst_out[21]), .B1(n1), .Y(
        n25) );
  INVX1 U124 ( .A(n26), .Y(n90) );
  AOI22X1 U125 ( .A0(inst_in[22]), .A1(n3), .B0(inst_out[22]), .B1(n1), .Y(n26) );
  INVX1 U126 ( .A(n27), .Y(n91) );
  AOI22X1 U127 ( .A0(inst_in[23]), .A1(n3), .B0(inst_out[23]), .B1(n1), .Y(n27) );
  INVX1 U128 ( .A(n28), .Y(n92) );
  AOI22X1 U129 ( .A0(inst_in[24]), .A1(n3), .B0(inst_out[24]), .B1(n1), .Y(n28) );
  INVX1 U130 ( .A(n29), .Y(n93) );
  AOI22X1 U131 ( .A0(inst_in[25]), .A1(n3), .B0(inst_out[25]), .B1(n1), .Y(n29) );
  INVX1 U132 ( .A(n33), .Y(n97) );
  AOI22X1 U133 ( .A0(inst_in[29]), .A1(n133), .B0(inst_out[29]), .B1(n1), .Y(
        n33) );
  INVX1 U134 ( .A(n36), .Y(n100) );
  AOI22X1 U135 ( .A0(pc_in[0]), .A1(n3), .B0(pc_out[0]), .B1(n1), .Y(n36) );
endmodule


module EXTENSION ( sign_ena, sel, imm_field, ext_out );
  input [2:0] sel;
  input [23:0] imm_field;
  output [31:0] ext_out;
  input sign_ena;
  wire   n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n43, n45, n46,
         n48, n50, n51, n52, n54, n56, n60, n61, n62, n63, n64, n66, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  assign ext_out[31] = ext_out[25];
  assign ext_out[30] = ext_out[25];
  assign ext_out[29] = ext_out[25];
  assign ext_out[28] = ext_out[25];
  assign ext_out[27] = ext_out[25];
  assign ext_out[26] = ext_out[25];

  NOR2X1 U2 ( .A(n50), .B(n62), .Y(n1) );
  NOR3X1 U3 ( .A(sel[0]), .B(sel[2]), .C(n66), .Y(n62) );
  BUFX3 U4 ( .A(n31), .Y(n2) );
  NOR2BX1 U5 ( .AN(n60), .B(sel[2]), .Y(n31) );
  INVX1 U6 ( .A(sel[2]), .Y(n45) );
  INVX1 U7 ( .A(n63), .Y(n40) );
  NAND3X1 U8 ( .A(n66), .B(n45), .C(sel[0]), .Y(n60) );
  INVX1 U9 ( .A(n54), .Y(n50) );
  NAND2X1 U10 ( .A(n64), .B(n63), .Y(n33) );
  INVX1 U11 ( .A(n51), .Y(n56) );
  NOR3X1 U12 ( .A(sel[1]), .B(sel[2]), .C(sel[0]), .Y(n63) );
  NAND3X1 U13 ( .A(sel[1]), .B(n45), .C(sel[0]), .Y(n54) );
  INVX1 U14 ( .A(sel[1]), .Y(n66) );
  OAI221XL U15 ( .A0(n1), .A1(n4), .B0(n2), .B1(n3), .C0(n33), .Y(ext_out[11])
         );
  OAI221XL U16 ( .A0(n1), .A1(n5), .B0(n2), .B1(n4), .C0(n33), .Y(ext_out[12])
         );
  OAI221XL U17 ( .A0(n1), .A1(n6), .B0(n2), .B1(n5), .C0(n33), .Y(ext_out[13])
         );
  NOR2X1 U18 ( .A(n46), .B(n7), .Y(n64) );
  INVX1 U19 ( .A(sign_ena), .Y(n46) );
  OAI31X1 U20 ( .A0(n45), .A1(n46), .A2(n13), .B0(n48), .Y(ext_out[25]) );
  OAI221XL U21 ( .A0(n54), .A1(n8), .B0(n7), .B1(n45), .C0(n56), .Y(
        ext_out[15]) );
  OAI221XL U22 ( .A0(n54), .A1(n9), .B0(n45), .B1(n8), .C0(n56), .Y(
        ext_out[16]) );
  OAI221XL U23 ( .A0(n54), .A1(n10), .B0(n45), .B1(n9), .C0(n56), .Y(
        ext_out[17]) );
  OAI221XL U24 ( .A0(n54), .A1(n11), .B0(n45), .B1(n10), .C0(n56), .Y(
        ext_out[18]) );
  OAI221XL U25 ( .A0(n54), .A1(n12), .B0(n45), .B1(n11), .C0(n56), .Y(
        ext_out[19]) );
  OAI221XL U26 ( .A0(n1), .A1(n7), .B0(n2), .B1(n6), .C0(n33), .Y(ext_out[14])
         );
  OAI21XL U27 ( .A0(n12), .A1(n45), .B0(n48), .Y(ext_out[20]) );
  OAI21XL U28 ( .A0(n13), .A1(n45), .B0(n48), .Y(ext_out[24]) );
  OAI31X1 U29 ( .A0(n60), .A1(n46), .A2(n6), .B0(n61), .Y(n51) );
  OAI21XL U30 ( .A0(n62), .A1(n63), .B0(n64), .Y(n61) );
  OAI222XL U31 ( .A0(n2), .A1(n52), .B0(n1), .B1(n43), .C0(n40), .C1(n4), .Y(
        ext_out[1]) );
  OAI222XL U32 ( .A0(n2), .A1(n43), .B0(n1), .B1(n41), .C0(n40), .C1(n5), .Y(
        ext_out[2]) );
  OAI222XL U33 ( .A0(n2), .A1(n41), .B0(n1), .B1(n38), .C0(n40), .C1(n6), .Y(
        ext_out[3]) );
  OAI22X1 U34 ( .A0(n40), .A1(n3), .B0(n1), .B1(n52), .Y(ext_out[0]) );
  OAI222XL U35 ( .A0(n2), .A1(n38), .B0(n1), .B1(n37), .C0(n7), .C1(n40), .Y(
        ext_out[4]) );
  OAI221XL U36 ( .A0(n1), .A1(n36), .B0(n2), .B1(n37), .C0(n33), .Y(ext_out[5]) );
  OAI221XL U37 ( .A0(n1), .A1(n35), .B0(n2), .B1(n36), .C0(n33), .Y(ext_out[6]) );
  OAI221XL U38 ( .A0(n1), .A1(n34), .B0(n2), .B1(n35), .C0(n33), .Y(ext_out[7]) );
  OAI221XL U39 ( .A0(n1), .A1(n32), .B0(n2), .B1(n34), .C0(n33), .Y(ext_out[8]) );
  OAI221XL U40 ( .A0(n1), .A1(n30), .B0(n2), .B1(n32), .C0(n33), .Y(ext_out[9]) );
  OAI221XL U41 ( .A0(n1), .A1(n3), .B0(n2), .B1(n30), .C0(n33), .Y(ext_out[10]) );
  INVX1 U42 ( .A(imm_field[14]), .Y(n7) );
  INVX1 U43 ( .A(imm_field[10]), .Y(n3) );
  INVX1 U44 ( .A(imm_field[13]), .Y(n6) );
  INVX1 U45 ( .A(imm_field[11]), .Y(n4) );
  INVX1 U46 ( .A(imm_field[12]), .Y(n5) );
  AOI31X1 U47 ( .A0(imm_field[19]), .A1(sign_ena), .A2(n50), .B0(n51), .Y(n48)
         );
  OAI2BB1X1 U48 ( .A0N(imm_field[20]), .A1N(sel[2]), .B0(n48), .Y(ext_out[21])
         );
  OAI2BB1X1 U49 ( .A0N(imm_field[21]), .A1N(sel[2]), .B0(n48), .Y(ext_out[22])
         );
  OAI2BB1X1 U50 ( .A0N(imm_field[22]), .A1N(sel[2]), .B0(n48), .Y(ext_out[23])
         );
  INVX1 U51 ( .A(imm_field[15]), .Y(n8) );
  INVX1 U52 ( .A(imm_field[16]), .Y(n9) );
  INVX1 U53 ( .A(imm_field[17]), .Y(n10) );
  INVX1 U54 ( .A(imm_field[18]), .Y(n11) );
  INVX1 U55 ( .A(imm_field[19]), .Y(n12) );
  INVX1 U56 ( .A(imm_field[23]), .Y(n13) );
  INVX1 U57 ( .A(imm_field[0]), .Y(n52) );
  INVX1 U58 ( .A(imm_field[1]), .Y(n43) );
  INVX1 U59 ( .A(imm_field[3]), .Y(n38) );
  INVX1 U60 ( .A(imm_field[2]), .Y(n41) );
  INVX1 U61 ( .A(imm_field[4]), .Y(n37) );
  INVX1 U62 ( .A(imm_field[5]), .Y(n36) );
  INVX1 U63 ( .A(imm_field[6]), .Y(n35) );
  INVX1 U64 ( .A(imm_field[7]), .Y(n34) );
  INVX1 U65 ( .A(imm_field[8]), .Y(n32) );
  INVX1 U66 ( .A(imm_field[9]), .Y(n30) );
endmodule


module CPU ( clk, rst );
  input clk, rst;
  wire   N29, stall, N33, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, sel_in2_out, sel_wb_reg2_out,
         sel_data1_in, branch_ena, sel_data2_in, reg_rw_in, sel_wb_in,
         data_rw_in, ena_data_in, sel_in2_in, ls_w_mode_in, reg_rw_in_control,
         sel_wb_in_control, data_rw_in_control, ena_data_in_control,
         sel_in2_in_control, ls_w_mode_in_control, compare, Jump_ena, flush,
         sel_alu_out, inst_out_31, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, sign_ena, reg_rw_reg2_out, sel_alu, ls_w_mode_out,
         ena_data_out, data_rw_out, sel_wb_out, reg_rw_out, ena_data_reg_out,
         data_rw_reg_out, sel_wb_reg_out, reg_rw_reg_out, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n176, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433;
  wire   [31:0] next_pc;
  wire   [31:0] source2;
  wire   [31:0] ext_reg_out;
  wire   [31:0] write_data;
  wire   [31:0] alu_result_reg_out;
  wire   [31:0] data_out_out;
  wire   [31:0] read_data1_out;
  wire   [1:0] forwardA;
  wire   [31:0] in1;
  wire   [31:0] alu_result_out;
  wire   [31:0] read_data2_out;
  wire   [1:0] forwardB;
  wire   [1:0] sel_data1;
  wire   [31:0] read_data1;
  wire   [31:0] result;
  wire   [1:0] sel_data3;
  wire   [31:0] read_data3_in;
  wire   [31:0] read_data3;
  wire   [31:0] read_data1_in;
  wire   [31:0] read_data2_in;
  wire   [31:0] read_data2;
  wire   [3:0] funct_in;
  wire   [3:0] funct_in_control;
  wire   [31:0] alu_result;
  wire   [31:0] data_in;
  wire   [31:0] read_data3_reg_out;
  wire   [9:5] inst_out;
  wire   [4:0] addr2;
  wire   [4:0] addr1;
  wire   [4:0] addr_dst;
  wire   [5:0] opcode;
  wire   [4:0] subopcode;
  wire   [31:0] pc_shift;
  wire   [31:0] next_pc_out;
  wire   [31:0] ext_out;
  wire   [2:0] sel;
  wire   [31:0] inst_in;
  wire   [4:0] addr_dst_reg2_out;
  wire   [3:0] funct_out;
  wire   [31:0] read_data3_out;
  wire   [4:0] addr_dst_out;
  wire   [4:0] addr1_out;
  wire   [4:0] addr2_out;
  wire   [31:0] inst_out2;
  wire   [4:0] addr_dst_reg_out;
  wire   [31:0] data_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29;

  EXTENSION ext ( .sign_ena(sign_ena), .sel(sel), .imm_field({addr_dst[3:0], 
        addr1, addr2[4], n431, n429, n427, n425, inst_out, subopcode}), 
        .ext_out(ext_out) );
  INST_MEM inst_mem ( .clk(clk), .pc({1'b0, 1'b0, next_pc[31:2]}), .inst_out(
        inst_in) );
  IFID ifid ( .pc_out(next_pc_out), .inst_out({inst_out_31, opcode, addr_dst, 
        addr1, addr2, inst_out, subopcode}), .pc_in(next_pc), .inst_in(inst_in), .clk(clk), .rst(rst), .flush(flush), .stall(stall) );
  REGISTER_FILE reg_file ( .clk(clk), .rst(rst), .reg_rw(reg_rw_reg2_out), 
        .reg_ena(1'b1), .addr1(addr1), .addr2({addr2[4], n431, n429, n427, 
        n425}), .addr_dst(addr_dst), .write_data(write_data), .write_addr(
        addr_dst_reg2_out), .read_data1(read_data1), .read_data2(read_data2), 
        .read_data3(read_data3) );
  CONTROLLER ctrl ( .funct(funct_in_control), .ls_w_mode(ls_w_mode_in_control), 
        .sign_ena(sign_ena), .sel_in2(sel_in2_in_control), .ena_data(
        ena_data_in_control), .data_rw(data_rw_in_control), .sel_wb(
        sel_wb_in_control), .reg_rw(reg_rw_in_control), .sel(sel), .opcode(
        opcode), .subopcode(subopcode), .read_data1(read_data1), .read_data2(
        read_data2), .clk(clk), .rst(rst), .sel_alu(sel_alu), .branch_ena(
        branch_ena), .Jump_ena(Jump_ena) );
  IDEX idex ( .ls_w_mode_out(ls_w_mode_out), .funct_out(funct_out), 
        .sel_in2_out(sel_in2_out), .ena_data_out(ena_data_out), .data_rw_out(
        data_rw_out), .sel_wb_out(sel_wb_out), .reg_rw_out(reg_rw_out), 
        .read_data1_out(read_data1_out), .read_data2_out(read_data2_out), 
        .read_data3_out(read_data3_out), .ext_out(ext_reg_out), .addr_dst_out(
        addr_dst_out), .ls_w_mode_in(ls_w_mode_in), .funct_in(funct_in), 
        .sel_in2_in(sel_in2_in), .ena_data_in(ena_data_in), .data_rw_in(
        data_rw_in), .sel_wb_in(sel_wb_in), .reg_rw_in(reg_rw_in), 
        .read_data1_in(read_data1_in), .read_data2_in(read_data2_in), 
        .addr_dst_in(addr_dst), .read_data3_in(read_data3_in), .ext_in(ext_out), .clk(clk), .rst(rst), .addr1_out(addr1_out), .addr1_in(addr1), .addr2_out(
        addr2_out), .addr2_in({addr2[4], n431, n429, n427, n425}), .inst_out({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, inst_out2[9:8], 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29}), .inst_in({
        inst_out_31, opcode, addr_dst, addr1, addr2[4], n431, n429, n427, n425, 
        inst_out, subopcode}), .sel_alu_out(sel_alu_out), .sel_alu_in(sel_alu)
         );
  ALU alu ( .ls_w_mode(ls_w_mode_out), .funct(funct_out), .sv(inst_out2[9:8]), 
        .source1(in1), .source2(source2), .alu_result(result) );
  EXMEM exmem ( .ena_data_out(ena_data_reg_out), .data_rw_out(data_rw_reg_out), 
        .sel_wb_out(sel_wb_reg_out), .reg_rw_out(reg_rw_reg_out), 
        .alu_result_out(alu_result_out), .read_data3_out(read_data3_reg_out), 
        .addr_dst_out(addr_dst_reg_out), .ena_data_in(ena_data_out), 
        .data_rw_in(data_rw_out), .sel_wb_in(sel_wb_out), .reg_rw_in(
        reg_rw_out), .alu_result_in(alu_result), .read_data3_in(read_data3_out), .addr_dst_in(addr_dst_out), .clk(clk), .rst(rst) );
  DATA_MEM data_mem ( .clk(clk), .rst(rst), .data_rw(data_rw_reg_out), 
        .ena_data(ena_data_reg_out), .addr(alu_result_out), .data_in(data_in), 
        .data_out(data_out) );
  MEMWB memwb ( .sel_wb_out(sel_wb_reg2_out), .reg_rw_out(reg_rw_reg2_out), 
        .addr_dst_out(addr_dst_reg2_out), .alu_result_out(alu_result_reg_out), 
        .data_out_out(data_out_out), .alu_result_in(alu_result_out), 
        .sel_wb_in(sel_wb_reg_out), .reg_rw_in(reg_rw_reg_out), .addr_dst_in(
        addr_dst_reg_out), .data_out_in(data_out), .clk(clk), .rst(rst) );
  Forward forwarding ( .forwardA(forwardA), .forwardB(forwardB), .addr2_out(
        addr2_out), .addr1_out(addr1_out), .addr_dst_reg_out(addr_dst_reg_out), 
        .addr_dst_reg2_out(addr_dst_reg2_out), .reg_rw_out_exe(reg_rw_reg_out), 
        .reg_rw_out_mem(reg_rw_reg2_out), .data_rw_reg_out(data_rw_reg_out), 
        .sel_data_in(N29), .addr_dst(addr_dst), .addr1(addr1), .branch_ena(
        branch_ena), .sel_data1(sel_data1), .sel_data3(sel_data3), 
        .addr_dst_out(addr_dst_out), .addr2({addr2[4], n431, n429, n427, n425}), .sel_data2_in(sel_data2_in), .sel_data1_in(sel_data1_in) );
  detection detect ( .stall(stall), .ena_data_out(ena_data_out), 
        .addr_dst_out(addr_dst_out), .addr1(addr1), .addr2({addr2[4], n431, 
        n429, n427, n425}) );
  CPU_DW01_add_0 add_216 ( .A(next_pc_out), .B(ext_out), .CI(1'b0), .SUM(
        pc_shift) );
  CPU_DW01_add_1 add_215 ( .A(next_pc), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N123, N122, N121, N120, N119, N118, 
        N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, 
        N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, 
        N92}) );
  CPU_DW01_cmp6_0 eq_218 ( .A(read_data3_in), .B(read_data1_in), .TC(1'b0), 
        .EQ(compare) );
  DFFRHQX1 \next_pc_reg[31]  ( .D(N66), .CK(clk), .RN(n72), .Q(next_pc[31]) );
  DFFRHQX1 \next_pc_reg[30]  ( .D(N65), .CK(clk), .RN(n72), .Q(next_pc[30]) );
  DFFRHQX1 \next_pc_reg[29]  ( .D(N64), .CK(clk), .RN(n72), .Q(next_pc[29]) );
  DFFRHQX1 \next_pc_reg[28]  ( .D(N63), .CK(clk), .RN(n72), .Q(next_pc[28]) );
  DFFRHQX1 \next_pc_reg[27]  ( .D(N62), .CK(clk), .RN(n72), .Q(next_pc[27]) );
  DFFRHQX1 \next_pc_reg[26]  ( .D(N61), .CK(clk), .RN(n72), .Q(next_pc[26]) );
  DFFRHQX1 \next_pc_reg[0]  ( .D(N35), .CK(clk), .RN(n72), .Q(next_pc[0]) );
  DFFRHQX1 \next_pc_reg[1]  ( .D(N36), .CK(clk), .RN(n72), .Q(next_pc[1]) );
  DFFRHQX1 \next_pc_reg[25]  ( .D(N60), .CK(clk), .RN(n72), .Q(next_pc[25]) );
  DFFRHQX1 \next_pc_reg[24]  ( .D(N59), .CK(clk), .RN(n72), .Q(next_pc[24]) );
  DFFRHQX1 \next_pc_reg[23]  ( .D(N58), .CK(clk), .RN(n72), .Q(next_pc[23]) );
  DFFRHQX1 \next_pc_reg[22]  ( .D(N57), .CK(clk), .RN(n72), .Q(next_pc[22]) );
  DFFRHQX1 \next_pc_reg[21]  ( .D(N56), .CK(clk), .RN(n72), .Q(next_pc[21]) );
  DFFRHQX1 \next_pc_reg[20]  ( .D(N55), .CK(clk), .RN(n72), .Q(next_pc[20]) );
  DFFRHQX1 \next_pc_reg[19]  ( .D(N54), .CK(clk), .RN(n72), .Q(next_pc[19]) );
  DFFRHQX1 \next_pc_reg[18]  ( .D(N53), .CK(clk), .RN(n72), .Q(next_pc[18]) );
  DFFRHQX1 \next_pc_reg[17]  ( .D(N52), .CK(clk), .RN(n72), .Q(next_pc[17]) );
  DFFRHQX1 \next_pc_reg[16]  ( .D(N51), .CK(clk), .RN(n72), .Q(next_pc[16]) );
  DFFRHQX1 \next_pc_reg[15]  ( .D(N50), .CK(clk), .RN(n72), .Q(next_pc[15]) );
  DFFRHQX1 \next_pc_reg[14]  ( .D(N49), .CK(clk), .RN(n72), .Q(next_pc[14]) );
  DFFRHQX1 \next_pc_reg[13]  ( .D(N48), .CK(clk), .RN(n72), .Q(next_pc[13]) );
  DFFRHQX1 \next_pc_reg[12]  ( .D(N47), .CK(clk), .RN(n72), .Q(next_pc[12]) );
  DFFRHQX1 \next_pc_reg[11]  ( .D(N46), .CK(clk), .RN(n72), .Q(next_pc[11]) );
  DFFRHQX1 \next_pc_reg[10]  ( .D(N45), .CK(clk), .RN(n72), .Q(next_pc[10]) );
  DFFRHQX1 \next_pc_reg[9]  ( .D(N44), .CK(clk), .RN(n72), .Q(next_pc[9]) );
  DFFRHQX1 \next_pc_reg[8]  ( .D(N43), .CK(clk), .RN(n72), .Q(next_pc[8]) );
  DFFRHQX1 \next_pc_reg[7]  ( .D(N42), .CK(clk), .RN(n72), .Q(next_pc[7]) );
  DFFRHQX1 \next_pc_reg[6]  ( .D(N41), .CK(clk), .RN(n72), .Q(next_pc[6]) );
  DFFRHQX1 \next_pc_reg[5]  ( .D(N40), .CK(clk), .RN(n72), .Q(next_pc[5]) );
  DFFRHQX1 \next_pc_reg[4]  ( .D(N39), .CK(clk), .RN(n72), .Q(next_pc[4]) );
  DFFRHQX1 \next_pc_reg[3]  ( .D(N38), .CK(clk), .RN(n72), .Q(next_pc[3]) );
  DFFRHQX1 \next_pc_reg[2]  ( .D(N37), .CK(clk), .RN(n72), .Q(next_pc[2]) );
  AND2X2 U120 ( .A(write_data[31]), .B(N29), .Y(n70) );
  AND2X2 U121 ( .A(read_data3_reg_out[31]), .B(n433), .Y(n71) );
  OR2X2 U122 ( .A(n70), .B(n71), .Y(data_in[31]) );
  AND2X2 U117 ( .A(write_data[30]), .B(N29), .Y(n68) );
  AND2X2 U118 ( .A(read_data3_reg_out[30]), .B(n433), .Y(n69) );
  OR2X2 U119 ( .A(n68), .B(n69), .Y(data_in[30]) );
  AND2X2 U114 ( .A(write_data[29]), .B(N29), .Y(n66) );
  AND2X2 U115 ( .A(read_data3_reg_out[29]), .B(n433), .Y(n67) );
  OR2X2 U116 ( .A(n66), .B(n67), .Y(data_in[29]) );
  AND2X2 U111 ( .A(write_data[28]), .B(N29), .Y(n64) );
  AND2X2 U112 ( .A(read_data3_reg_out[28]), .B(n433), .Y(n65) );
  OR2X2 U113 ( .A(n64), .B(n65), .Y(data_in[28]) );
  AND2X2 U108 ( .A(write_data[27]), .B(N29), .Y(n62) );
  AND2X2 U109 ( .A(read_data3_reg_out[27]), .B(n433), .Y(n63) );
  OR2X2 U110 ( .A(n62), .B(n63), .Y(data_in[27]) );
  AND2X2 U105 ( .A(write_data[26]), .B(N29), .Y(n60) );
  AND2X2 U106 ( .A(read_data3_reg_out[26]), .B(n433), .Y(n61) );
  OR2X2 U107 ( .A(n60), .B(n61), .Y(data_in[26]) );
  AND2X2 U102 ( .A(write_data[25]), .B(N29), .Y(n58) );
  AND2X2 U103 ( .A(read_data3_reg_out[25]), .B(n433), .Y(n59) );
  OR2X2 U104 ( .A(n58), .B(n59), .Y(data_in[25]) );
  AND2X2 U99 ( .A(write_data[24]), .B(N29), .Y(n56) );
  AND2X2 U100 ( .A(read_data3_reg_out[24]), .B(n433), .Y(n57) );
  OR2X2 U101 ( .A(n56), .B(n57), .Y(data_in[24]) );
  AND2X2 U96 ( .A(write_data[23]), .B(N29), .Y(n54) );
  AND2X2 U97 ( .A(read_data3_reg_out[23]), .B(n433), .Y(n55) );
  OR2X2 U98 ( .A(n54), .B(n55), .Y(data_in[23]) );
  AND2X2 U93 ( .A(write_data[22]), .B(N29), .Y(n52) );
  AND2X2 U94 ( .A(read_data3_reg_out[22]), .B(n433), .Y(n53) );
  OR2X2 U95 ( .A(n52), .B(n53), .Y(data_in[22]) );
  AND2X2 U90 ( .A(write_data[21]), .B(N29), .Y(n50) );
  AND2X2 U91 ( .A(read_data3_reg_out[21]), .B(n433), .Y(n51) );
  OR2X2 U92 ( .A(n50), .B(n51), .Y(data_in[21]) );
  AND2X2 U87 ( .A(write_data[20]), .B(N29), .Y(n48) );
  AND2X2 U88 ( .A(read_data3_reg_out[20]), .B(n433), .Y(n49) );
  OR2X2 U89 ( .A(n48), .B(n49), .Y(data_in[20]) );
  AND2X2 U84 ( .A(write_data[19]), .B(N29), .Y(n46) );
  AND2X2 U85 ( .A(read_data3_reg_out[19]), .B(n433), .Y(n47) );
  OR2X2 U86 ( .A(n46), .B(n47), .Y(data_in[19]) );
  AND2X2 U81 ( .A(write_data[18]), .B(N29), .Y(n44) );
  AND2X2 U82 ( .A(read_data3_reg_out[18]), .B(n433), .Y(n45) );
  OR2X2 U83 ( .A(n44), .B(n45), .Y(data_in[18]) );
  AND2X2 U78 ( .A(write_data[17]), .B(N29), .Y(n42) );
  AND2X2 U79 ( .A(read_data3_reg_out[17]), .B(n433), .Y(n43) );
  OR2X2 U80 ( .A(n42), .B(n43), .Y(data_in[17]) );
  AND2X2 U75 ( .A(write_data[16]), .B(N29), .Y(n40) );
  AND2X2 U76 ( .A(read_data3_reg_out[16]), .B(n433), .Y(n41) );
  OR2X2 U77 ( .A(n40), .B(n41), .Y(data_in[16]) );
  AND2X2 U72 ( .A(write_data[15]), .B(N29), .Y(n38) );
  AND2X2 U73 ( .A(read_data3_reg_out[15]), .B(n433), .Y(n39) );
  OR2X2 U74 ( .A(n38), .B(n39), .Y(data_in[15]) );
  AND2X2 U69 ( .A(write_data[14]), .B(N29), .Y(n36) );
  AND2X2 U70 ( .A(read_data3_reg_out[14]), .B(n433), .Y(n37) );
  OR2X2 U71 ( .A(n36), .B(n37), .Y(data_in[14]) );
  AND2X2 U66 ( .A(write_data[13]), .B(N29), .Y(n34) );
  AND2X2 U67 ( .A(read_data3_reg_out[13]), .B(n433), .Y(n35) );
  OR2X2 U68 ( .A(n34), .B(n35), .Y(data_in[13]) );
  AND2X2 U63 ( .A(write_data[12]), .B(N29), .Y(n32) );
  AND2X2 U64 ( .A(read_data3_reg_out[12]), .B(n433), .Y(n33) );
  OR2X2 U65 ( .A(n32), .B(n33), .Y(data_in[12]) );
  AND2X2 U60 ( .A(write_data[11]), .B(N29), .Y(n30) );
  AND2X2 U61 ( .A(read_data3_reg_out[11]), .B(n433), .Y(n31) );
  OR2X2 U62 ( .A(n30), .B(n31), .Y(data_in[11]) );
  AND2X2 U57 ( .A(write_data[10]), .B(N29), .Y(n28) );
  AND2X2 U58 ( .A(read_data3_reg_out[10]), .B(n433), .Y(n29) );
  OR2X2 U59 ( .A(n28), .B(n29), .Y(data_in[10]) );
  AND2X2 U54 ( .A(write_data[9]), .B(N29), .Y(n26) );
  AND2X2 U55 ( .A(read_data3_reg_out[9]), .B(n433), .Y(n27) );
  OR2X2 U56 ( .A(n26), .B(n27), .Y(data_in[9]) );
  AND2X2 U51 ( .A(write_data[8]), .B(N29), .Y(n24) );
  AND2X2 U52 ( .A(read_data3_reg_out[8]), .B(n433), .Y(n25) );
  OR2X2 U53 ( .A(n24), .B(n25), .Y(data_in[8]) );
  AND2X2 U48 ( .A(write_data[7]), .B(N29), .Y(n22) );
  AND2X2 U49 ( .A(read_data3_reg_out[7]), .B(n433), .Y(n23) );
  OR2X2 U50 ( .A(n22), .B(n23), .Y(data_in[7]) );
  AND2X2 U45 ( .A(write_data[6]), .B(N29), .Y(n20) );
  AND2X2 U46 ( .A(read_data3_reg_out[6]), .B(n433), .Y(n21) );
  OR2X2 U47 ( .A(n20), .B(n21), .Y(data_in[6]) );
  AND2X2 U42 ( .A(write_data[5]), .B(N29), .Y(n18) );
  AND2X2 U43 ( .A(read_data3_reg_out[5]), .B(n433), .Y(n19) );
  OR2X2 U44 ( .A(n18), .B(n19), .Y(data_in[5]) );
  AND2X2 U39 ( .A(write_data[4]), .B(N29), .Y(n16) );
  AND2X2 U40 ( .A(read_data3_reg_out[4]), .B(n433), .Y(n17) );
  OR2X2 U41 ( .A(n16), .B(n17), .Y(data_in[4]) );
  AND2X2 U36 ( .A(write_data[3]), .B(N29), .Y(n14) );
  AND2X2 U37 ( .A(read_data3_reg_out[3]), .B(n433), .Y(n15) );
  OR2X2 U38 ( .A(n14), .B(n15), .Y(data_in[3]) );
  AND2X2 U33 ( .A(write_data[2]), .B(N29), .Y(n12) );
  AND2X2 U34 ( .A(read_data3_reg_out[2]), .B(n433), .Y(n13) );
  OR2X2 U35 ( .A(n12), .B(n13), .Y(data_in[2]) );
  AND2X2 U30 ( .A(write_data[1]), .B(N29), .Y(n10) );
  AND2X2 U31 ( .A(read_data3_reg_out[1]), .B(n433), .Y(n11) );
  OR2X2 U32 ( .A(n10), .B(n11), .Y(data_in[1]) );
  AND2X2 U27 ( .A(write_data[0]), .B(N29), .Y(n8) );
  AND2X2 U28 ( .A(read_data3_reg_out[0]), .B(n433), .Y(n9) );
  OR2X2 U29 ( .A(n8), .B(n9), .Y(data_in[0]) );
  AND2X2 U652 ( .A(n172), .B(n424), .Y(n353) );
  NOR2X1 U653 ( .A(n210), .B(sel_data3[1]), .Y(n354) );
  NOR2X1 U654 ( .A(sel_data3[0]), .B(sel_data3[1]), .Y(n355) );
  NAND2X1 U655 ( .A(sel_data3[1]), .B(sel_data3[0]), .Y(n356) );
  NAND2X1 U656 ( .A(sel_data3[1]), .B(n210), .Y(n357) );
  INVX1 U657 ( .A(n362), .Y(n364) );
  INVX1 U658 ( .A(n362), .Y(n365) );
  INVX1 U659 ( .A(n362), .Y(n363) );
  INVX1 U660 ( .A(n360), .Y(n361) );
  INVX1 U661 ( .A(n366), .Y(n367) );
  INVX1 U662 ( .A(n375), .Y(n376) );
  INVX1 U663 ( .A(n371), .Y(n373) );
  INVX1 U664 ( .A(n371), .Y(n374) );
  INVX1 U665 ( .A(n371), .Y(n372) );
  INVX1 U666 ( .A(n377), .Y(n378) );
  INVX1 U667 ( .A(n366), .Y(n368) );
  INVX1 U668 ( .A(n370), .Y(n375) );
  INVX1 U669 ( .A(n369), .Y(n371) );
  INVX1 U670 ( .A(n359), .Y(n362) );
  INVX1 U671 ( .A(n358), .Y(n360) );
  INVX1 U672 ( .A(n320), .Y(n377) );
  INVX1 U673 ( .A(n319), .Y(n366) );
  INVX1 U674 ( .A(n382), .Y(n383) );
  INVX1 U675 ( .A(n381), .Y(n384) );
  INVX1 U676 ( .A(n381), .Y(n385) );
  INVX1 U677 ( .A(n381), .Y(n386) );
  INVX1 U678 ( .A(n382), .Y(n387) );
  INVX1 U679 ( .A(n382), .Y(n388) );
  NOR2X1 U680 ( .A(n352), .B(stall), .Y(n320) );
  INVX1 U681 ( .A(n283), .Y(n381) );
  INVX1 U682 ( .A(n283), .Y(n382) );
  NOR2X1 U683 ( .A(flush), .B(stall), .Y(n319) );
  INVX1 U684 ( .A(n352), .Y(flush) );
  NOR2X1 U685 ( .A(n352), .B(stall), .Y(n370) );
  NOR2X1 U686 ( .A(n352), .B(stall), .Y(n369) );
  NOR2X1 U687 ( .A(flush), .B(stall), .Y(n359) );
  NOR2X1 U688 ( .A(flush), .B(stall), .Y(n358) );
  BUFX3 U689 ( .A(n285), .Y(n390) );
  BUFX3 U690 ( .A(n285), .Y(n389) );
  INVX1 U691 ( .A(n74), .Y(n402) );
  INVX1 U692 ( .A(n74), .Y(n401) );
  INVX1 U693 ( .A(n74), .Y(n400) );
  INVX1 U694 ( .A(n423), .Y(n414) );
  INVX1 U695 ( .A(n423), .Y(n415) );
  INVX1 U696 ( .A(result[28]), .Y(n238) );
  INVX1 U697 ( .A(result[26]), .Y(n242) );
  INVX1 U698 ( .A(result[27]), .Y(n240) );
  INVX1 U699 ( .A(result[22]), .Y(n250) );
  INVX1 U700 ( .A(result[25]), .Y(n244) );
  INVX1 U701 ( .A(result[29]), .Y(n236) );
  INVX1 U702 ( .A(result[24]), .Y(n246) );
  INVX1 U703 ( .A(result[30]), .Y(n232) );
  INVX1 U704 ( .A(result[23]), .Y(n248) );
  INVX1 U705 ( .A(result[21]), .Y(n252) );
  INVX1 U706 ( .A(result[31]), .Y(n230) );
  INVX1 U707 ( .A(n423), .Y(n416) );
  INVX1 U708 ( .A(n410), .Y(n422) );
  INVX1 U709 ( .A(n410), .Y(n421) );
  INVX1 U710 ( .A(n409), .Y(n419) );
  INVX1 U711 ( .A(n409), .Y(n417) );
  INVX1 U712 ( .A(n409), .Y(n418) );
  INVX1 U713 ( .A(result[9]), .Y(n213) );
  INVX1 U714 ( .A(result[8]), .Y(n218) );
  INVX1 U715 ( .A(result[7]), .Y(n220) );
  INVX1 U716 ( .A(result[6]), .Y(n222) );
  INVX1 U717 ( .A(result[10]), .Y(n276) );
  INVX1 U718 ( .A(result[16]), .Y(n264) );
  INVX1 U719 ( .A(result[18]), .Y(n260) );
  INVX1 U720 ( .A(result[12]), .Y(n272) );
  INVX1 U721 ( .A(result[13]), .Y(n270) );
  INVX1 U722 ( .A(result[19]), .Y(n258) );
  INVX1 U723 ( .A(result[20]), .Y(n254) );
  INVX1 U724 ( .A(result[11]), .Y(n274) );
  INVX1 U725 ( .A(result[17]), .Y(n262) );
  INVX1 U726 ( .A(result[15]), .Y(n266) );
  INVX1 U727 ( .A(result[14]), .Y(n268) );
  INVX1 U728 ( .A(result[0]), .Y(n278) );
  INVX1 U729 ( .A(result[1]), .Y(n256) );
  INVX1 U730 ( .A(result[2]), .Y(n234) );
  INVX1 U731 ( .A(result[3]), .Y(n228) );
  INVX1 U732 ( .A(result[4]), .Y(n226) );
  INVX1 U733 ( .A(result[5]), .Y(n224) );
  INVX1 U734 ( .A(n409), .Y(n420) );
  INVX1 U735 ( .A(sel_data3[0]), .Y(n210) );
  BUFX3 U736 ( .A(n216), .Y(n394) );
  BUFX3 U737 ( .A(n216), .Y(n393) );
  NOR2BX1 U738 ( .AN(reg_rw_in_control), .B(stall), .Y(reg_rw_in) );
  NOR2BX1 U739 ( .AN(sel_wb_in_control), .B(stall), .Y(sel_wb_in) );
  NOR2BX1 U740 ( .AN(ena_data_in_control), .B(stall), .Y(ena_data_in) );
  NOR2BX1 U741 ( .AN(ls_w_mode_in_control), .B(stall), .Y(ls_w_mode_in) );
  AOI21X1 U742 ( .A0(compare), .A1(branch_ena), .B0(Jump_ena), .Y(n352) );
  NAND3BX1 U743 ( .AN(forwardB[0]), .B(n424), .C(forwardB[1]), .Y(n74) );
  BUFX3 U744 ( .A(n282), .Y(n380) );
  NAND2BX1 U745 ( .AN(forwardA[0]), .B(forwardA[1]), .Y(n282) );
  NAND2BX1 U746 ( .AN(forwardA[1]), .B(forwardA[0]), .Y(n283) );
  XNOR2X1 U747 ( .A(forwardA[0]), .B(forwardA[1]), .Y(n285) );
  BUFX3 U748 ( .A(n75), .Y(n408) );
  NAND3BX1 U749 ( .AN(forwardB[1]), .B(n424), .C(forwardB[0]), .Y(n75) );
  XNOR2X1 U750 ( .A(forwardB[0]), .B(forwardB[1]), .Y(n172) );
  INVX1 U751 ( .A(n411), .Y(n423) );
  INVX1 U752 ( .A(n412), .Y(n411) );
  INVX1 U753 ( .A(n412), .Y(n410) );
  INVX1 U754 ( .A(n413), .Y(n409) );
  BUFX3 U755 ( .A(n212), .Y(n391) );
  NAND3BX1 U756 ( .AN(sel_data1[0]), .B(branch_ena), .C(sel_data1[1]), .Y(n212) );
  BUFX3 U757 ( .A(n214), .Y(n392) );
  NAND3BX1 U758 ( .AN(sel_data1[1]), .B(branch_ena), .C(sel_data1[0]), .Y(n214) );
  INVX1 U759 ( .A(n281), .Y(n216) );
  AOI32X1 U760 ( .A0(sel_data1[0]), .A1(branch_ena), .A2(sel_data1[1]), .B0(
        n280), .B1(sel_data1_in), .Y(n281) );
  INVX1 U761 ( .A(n169), .Y(write_data[0]) );
  INVX1 U762 ( .A(n136), .Y(write_data[1]) );
  INVX1 U763 ( .A(n103), .Y(write_data[2]) );
  INVX1 U764 ( .A(n94), .Y(write_data[3]) );
  INVX1 U765 ( .A(n88), .Y(write_data[5]) );
  INVX1 U766 ( .A(n85), .Y(write_data[6]) );
  INVX1 U767 ( .A(n82), .Y(write_data[7]) );
  INVX1 U768 ( .A(n79), .Y(write_data[8]) );
  INVX1 U769 ( .A(n73), .Y(write_data[9]) );
  INVX1 U770 ( .A(n166), .Y(write_data[10]) );
  INVX1 U771 ( .A(n163), .Y(write_data[11]) );
  INVX1 U772 ( .A(n160), .Y(write_data[12]) );
  INVX1 U773 ( .A(n157), .Y(write_data[13]) );
  INVX1 U774 ( .A(n154), .Y(write_data[14]) );
  INVX1 U775 ( .A(n151), .Y(write_data[15]) );
  INVX1 U776 ( .A(n148), .Y(write_data[16]) );
  INVX1 U777 ( .A(n145), .Y(write_data[17]) );
  INVX1 U778 ( .A(n142), .Y(write_data[18]) );
  INVX1 U779 ( .A(n139), .Y(write_data[19]) );
  INVX1 U780 ( .A(n133), .Y(write_data[20]) );
  INVX1 U781 ( .A(n130), .Y(write_data[21]) );
  INVX1 U782 ( .A(n127), .Y(write_data[22]) );
  INVX1 U783 ( .A(n124), .Y(write_data[23]) );
  INVX1 U784 ( .A(n121), .Y(write_data[24]) );
  INVX1 U785 ( .A(n118), .Y(write_data[25]) );
  INVX1 U786 ( .A(n115), .Y(write_data[26]) );
  INVX1 U787 ( .A(n112), .Y(write_data[27]) );
  INVX1 U788 ( .A(n109), .Y(write_data[28]) );
  INVX1 U789 ( .A(n106), .Y(write_data[29]) );
  INVX1 U790 ( .A(n100), .Y(write_data[30]) );
  INVX1 U791 ( .A(n97), .Y(write_data[31]) );
  OAI32X1 U792 ( .A0(n280), .A1(sel_data1[1]), .A2(sel_data1[0]), .B0(
        sel_data1_in), .B1(branch_ena), .Y(n396) );
  OAI32X1 U793 ( .A0(n280), .A1(sel_data1[1]), .A2(sel_data1[0]), .B0(
        sel_data1_in), .B1(branch_ena), .Y(n217) );
  OAI32X1 U794 ( .A0(n280), .A1(sel_data1[1]), .A2(sel_data1[0]), .B0(
        sel_data1_in), .B1(branch_ena), .Y(n395) );
  INVX1 U795 ( .A(branch_ena), .Y(n280) );
  BUFX3 U796 ( .A(n211), .Y(n398) );
  BUFX3 U797 ( .A(n211), .Y(n399) );
  INVX1 U798 ( .A(n91), .Y(write_data[4]) );
  NOR2BX1 U799 ( .AN(data_rw_in_control), .B(stall), .Y(data_rw_in) );
  NOR2BX1 U800 ( .AN(sel_in2_in_control), .B(stall), .Y(sel_in2_in) );
  NOR2BX1 U801 ( .AN(funct_in_control[0]), .B(stall), .Y(funct_in[0]) );
  NOR2BX1 U802 ( .AN(funct_in_control[1]), .B(stall), .Y(funct_in[1]) );
  BUFX3 U803 ( .A(n211), .Y(n397) );
  INVX1 U804 ( .A(N29), .Y(n433) );
  OAI221XL U805 ( .A0(n79), .A1(n406), .B0(n408), .B1(n80), .C0(n81), .Y(
        source2[8]) );
  AOI22X1 U806 ( .A0(read_data2_out[8]), .A1(n353), .B0(ext_reg_out[8]), .B1(
        sel_in2_out), .Y(n81) );
  OAI221XL U807 ( .A0(n82), .A1(n405), .B0(n408), .B1(n83), .C0(n84), .Y(
        source2[7]) );
  AOI22X1 U808 ( .A0(read_data2_out[7]), .A1(n353), .B0(ext_reg_out[7]), .B1(
        sel_in2_out), .Y(n84) );
  OAI221XL U809 ( .A0(n85), .A1(n406), .B0(n408), .B1(n86), .C0(n87), .Y(
        source2[6]) );
  AOI22X1 U810 ( .A0(read_data2_out[6]), .A1(n353), .B0(ext_reg_out[6]), .B1(
        sel_in2_out), .Y(n87) );
  OAI221XL U811 ( .A0(n166), .A1(n404), .B0(n408), .B1(n167), .C0(n168), .Y(
        source2[10]) );
  AOI22X1 U812 ( .A0(read_data2_out[10]), .A1(n353), .B0(ext_reg_out[10]), 
        .B1(sel_in2_out), .Y(n168) );
  AOI22X1 U813 ( .A0(alu_result_reg_out[0]), .A1(n414), .B0(data_out_out[0]), 
        .B1(n422), .Y(n169) );
  AOI22X1 U814 ( .A0(alu_result_reg_out[1]), .A1(n414), .B0(data_out_out[1]), 
        .B1(n421), .Y(n136) );
  AOI22X1 U815 ( .A0(alu_result_reg_out[2]), .A1(n415), .B0(data_out_out[2]), 
        .B1(n419), .Y(n103) );
  AOI22X1 U816 ( .A0(alu_result_reg_out[3]), .A1(n416), .B0(data_out_out[3]), 
        .B1(n418), .Y(n94) );
  AOI22X1 U817 ( .A0(alu_result_reg_out[4]), .A1(n416), .B0(data_out_out[4]), 
        .B1(n417), .Y(n91) );
  AOI22X1 U818 ( .A0(alu_result_reg_out[5]), .A1(n416), .B0(data_out_out[5]), 
        .B1(n417), .Y(n88) );
  AOI22X1 U819 ( .A0(alu_result_reg_out[6]), .A1(n416), .B0(data_out_out[6]), 
        .B1(n420), .Y(n85) );
  AOI22X1 U820 ( .A0(alu_result_reg_out[7]), .A1(n416), .B0(data_out_out[7]), 
        .B1(n420), .Y(n82) );
  AOI22X1 U821 ( .A0(alu_result_reg_out[8]), .A1(n416), .B0(data_out_out[8]), 
        .B1(n420), .Y(n79) );
  OAI221XL U822 ( .A0(n130), .A1(n356), .B0(n131), .B1(n357), .C0(n196), .Y(
        read_data3_in[21]) );
  AOI22X1 U823 ( .A0(result[21]), .A1(n354), .B0(read_data3[21]), .B1(n355), 
        .Y(n196) );
  OAI221XL U824 ( .A0(n127), .A1(n356), .B0(n128), .B1(n357), .C0(n195), .Y(
        read_data3_in[22]) );
  AOI22X1 U825 ( .A0(result[22]), .A1(n354), .B0(read_data3[22]), .B1(n355), 
        .Y(n195) );
  OAI221XL U826 ( .A0(n124), .A1(n356), .B0(n125), .B1(n357), .C0(n194), .Y(
        read_data3_in[23]) );
  AOI22X1 U827 ( .A0(result[23]), .A1(n354), .B0(read_data3[23]), .B1(n355), 
        .Y(n194) );
  OAI221XL U828 ( .A0(n121), .A1(n356), .B0(n122), .B1(n357), .C0(n193), .Y(
        read_data3_in[24]) );
  AOI22X1 U829 ( .A0(result[24]), .A1(n354), .B0(read_data3[24]), .B1(n355), 
        .Y(n193) );
  OAI221XL U830 ( .A0(n118), .A1(n356), .B0(n119), .B1(n357), .C0(n192), .Y(
        read_data3_in[25]) );
  AOI22X1 U831 ( .A0(result[25]), .A1(n354), .B0(read_data3[25]), .B1(n355), 
        .Y(n192) );
  OAI221XL U832 ( .A0(n115), .A1(n356), .B0(n116), .B1(n357), .C0(n191), .Y(
        read_data3_in[26]) );
  AOI22X1 U833 ( .A0(result[26]), .A1(n354), .B0(read_data3[26]), .B1(n355), 
        .Y(n191) );
  OAI221XL U834 ( .A0(n112), .A1(n356), .B0(n113), .B1(n357), .C0(n190), .Y(
        read_data3_in[27]) );
  AOI22X1 U835 ( .A0(result[27]), .A1(n354), .B0(read_data3[27]), .B1(n355), 
        .Y(n190) );
  OAI221XL U836 ( .A0(n109), .A1(n356), .B0(n110), .B1(n357), .C0(n189), .Y(
        read_data3_in[28]) );
  AOI22X1 U837 ( .A0(result[28]), .A1(n354), .B0(read_data3[28]), .B1(n355), 
        .Y(n189) );
  OAI221XL U838 ( .A0(n106), .A1(n356), .B0(n107), .B1(n357), .C0(n188), .Y(
        read_data3_in[29]) );
  AOI22X1 U839 ( .A0(result[29]), .A1(n354), .B0(read_data3[29]), .B1(n355), 
        .Y(n188) );
  OAI221XL U840 ( .A0(n100), .A1(n356), .B0(n101), .B1(n357), .C0(n186), .Y(
        read_data3_in[30]) );
  AOI22X1 U841 ( .A0(result[30]), .A1(n354), .B0(read_data3[30]), .B1(n355), 
        .Y(n186) );
  OAI221XL U842 ( .A0(n97), .A1(n356), .B0(n98), .B1(n357), .C0(n185), .Y(
        read_data3_in[31]) );
  AOI22X1 U843 ( .A0(result[31]), .A1(n354), .B0(read_data3[31]), .B1(n355), 
        .Y(n185) );
  OAI221XL U844 ( .A0(n131), .A1(n391), .B0(n252), .B1(n392), .C0(n253), .Y(
        read_data1_in[21]) );
  AOI22X1 U845 ( .A0(n394), .A1(write_data[21]), .B0(read_data1[21]), .B1(n217), .Y(n253) );
  OAI221XL U846 ( .A0(n128), .A1(n391), .B0(n250), .B1(n392), .C0(n251), .Y(
        read_data1_in[22]) );
  AOI22X1 U847 ( .A0(n394), .A1(write_data[22]), .B0(read_data1[22]), .B1(n396), .Y(n251) );
  OAI221XL U848 ( .A0(n125), .A1(n391), .B0(n248), .B1(n392), .C0(n249), .Y(
        read_data1_in[23]) );
  AOI22X1 U849 ( .A0(n393), .A1(write_data[23]), .B0(read_data1[23]), .B1(n396), .Y(n249) );
  OAI221XL U850 ( .A0(n122), .A1(n391), .B0(n246), .B1(n392), .C0(n247), .Y(
        read_data1_in[24]) );
  AOI22X1 U851 ( .A0(n393), .A1(write_data[24]), .B0(read_data1[24]), .B1(n217), .Y(n247) );
  OAI221XL U852 ( .A0(n119), .A1(n391), .B0(n244), .B1(n392), .C0(n245), .Y(
        read_data1_in[25]) );
  AOI22X1 U853 ( .A0(n393), .A1(write_data[25]), .B0(read_data1[25]), .B1(n217), .Y(n245) );
  OAI221XL U854 ( .A0(n116), .A1(n391), .B0(n242), .B1(n392), .C0(n243), .Y(
        read_data1_in[26]) );
  AOI22X1 U855 ( .A0(n393), .A1(write_data[26]), .B0(read_data1[26]), .B1(n217), .Y(n243) );
  OAI221XL U856 ( .A0(n113), .A1(n391), .B0(n240), .B1(n392), .C0(n241), .Y(
        read_data1_in[27]) );
  AOI22X1 U857 ( .A0(n393), .A1(write_data[27]), .B0(read_data1[27]), .B1(n217), .Y(n241) );
  OAI221XL U858 ( .A0(n110), .A1(n391), .B0(n238), .B1(n392), .C0(n239), .Y(
        read_data1_in[28]) );
  AOI22X1 U859 ( .A0(n393), .A1(write_data[28]), .B0(read_data1[28]), .B1(n217), .Y(n239) );
  OAI221XL U860 ( .A0(n107), .A1(n391), .B0(n236), .B1(n392), .C0(n237), .Y(
        read_data1_in[29]) );
  AOI22X1 U861 ( .A0(n393), .A1(write_data[29]), .B0(read_data1[29]), .B1(n217), .Y(n237) );
  OAI221XL U862 ( .A0(n101), .A1(n391), .B0(n232), .B1(n392), .C0(n233), .Y(
        read_data1_in[30]) );
  AOI22X1 U863 ( .A0(n393), .A1(write_data[30]), .B0(read_data1[30]), .B1(n395), .Y(n233) );
  OAI221XL U864 ( .A0(n98), .A1(n391), .B0(n230), .B1(n392), .C0(n231), .Y(
        read_data1_in[31]) );
  AOI22X1 U865 ( .A0(n393), .A1(write_data[31]), .B0(read_data1[31]), .B1(n395), .Y(n231) );
  OAI2BB1X1 U866 ( .A0N(next_pc[18]), .A1N(stall), .B0(n333), .Y(N53) );
  AOI22X1 U867 ( .A0(N110), .A1(n367), .B0(pc_shift[18]), .B1(n379), .Y(n333)
         );
  OAI2BB1X1 U868 ( .A0N(next_pc[19]), .A1N(stall), .B0(n332), .Y(N54) );
  AOI22X1 U869 ( .A0(N111), .A1(n368), .B0(pc_shift[19]), .B1(n379), .Y(n332)
         );
  INVX1 U870 ( .A(n377), .Y(n379) );
  OAI2BB1X1 U871 ( .A0N(next_pc[20]), .A1N(stall), .B0(n331), .Y(N55) );
  AOI22X1 U872 ( .A0(N112), .A1(n368), .B0(pc_shift[20]), .B1(n379), .Y(n331)
         );
  OAI2BB1X1 U873 ( .A0N(next_pc[21]), .A1N(stall), .B0(n330), .Y(N56) );
  AOI22X1 U874 ( .A0(N113), .A1(n368), .B0(pc_shift[21]), .B1(n379), .Y(n330)
         );
  OAI221XL U875 ( .A0(n73), .A1(n406), .B0(n408), .B1(n76), .C0(n77), .Y(
        source2[9]) );
  AOI22X1 U876 ( .A0(read_data2_out[9]), .A1(n353), .B0(sel_in2_out), .B1(
        ext_reg_out[9]), .Y(n77) );
  OAI221XL U877 ( .A0(n91), .A1(n405), .B0(n408), .B1(n92), .C0(n93), .Y(
        source2[4]) );
  AOI22X1 U878 ( .A0(read_data2_out[4]), .A1(n353), .B0(ext_reg_out[4]), .B1(
        sel_in2_out), .Y(n93) );
  OAI221XL U879 ( .A0(n103), .A1(n403), .B0(n408), .B1(n104), .C0(n105), .Y(
        source2[2]) );
  AOI22X1 U880 ( .A0(read_data2_out[2]), .A1(n353), .B0(ext_reg_out[2]), .B1(
        sel_in2_out), .Y(n105) );
  OAI221XL U881 ( .A0(n94), .A1(n405), .B0(n408), .B1(n95), .C0(n96), .Y(
        source2[3]) );
  AOI22X1 U882 ( .A0(read_data2_out[3]), .A1(n353), .B0(ext_reg_out[3]), .B1(
        sel_in2_out), .Y(n96) );
  INVX1 U883 ( .A(alu_result_out[0]), .Y(n170) );
  INVX1 U884 ( .A(alu_result_out[1]), .Y(n137) );
  INVX1 U885 ( .A(alu_result_out[2]), .Y(n104) );
  OAI221XL U886 ( .A0(n94), .A1(n380), .B0(n95), .B1(n384), .C0(n292), .Y(
        in1[3]) );
  NAND2X1 U887 ( .A(read_data1_out[3]), .B(n390), .Y(n292) );
  OAI221XL U888 ( .A0(n91), .A1(n380), .B0(n92), .B1(n385), .C0(n291), .Y(
        in1[4]) );
  NAND2X1 U889 ( .A(read_data1_out[4]), .B(n389), .Y(n291) );
  OAI221XL U890 ( .A0(n88), .A1(n380), .B0(n89), .B1(n386), .C0(n290), .Y(
        in1[5]) );
  NAND2X1 U891 ( .A(read_data1_out[5]), .B(n390), .Y(n290) );
  OAI221XL U892 ( .A0(n85), .A1(n380), .B0(n86), .B1(n387), .C0(n289), .Y(
        in1[6]) );
  NAND2X1 U893 ( .A(read_data1_out[6]), .B(n389), .Y(n289) );
  OAI221XL U894 ( .A0(n82), .A1(n380), .B0(n83), .B1(n387), .C0(n288), .Y(
        in1[7]) );
  NAND2X1 U895 ( .A(read_data1_out[7]), .B(n390), .Y(n288) );
  OAI221XL U896 ( .A0(n79), .A1(n380), .B0(n80), .B1(n387), .C0(n287), .Y(
        in1[8]) );
  NAND2X1 U897 ( .A(read_data1_out[8]), .B(n389), .Y(n287) );
  OAI221XL U898 ( .A0(n73), .A1(n380), .B0(n76), .B1(n387), .C0(n284), .Y(
        in1[9]) );
  NAND2X1 U899 ( .A(read_data1_out[9]), .B(n390), .Y(n284) );
  OAI221XL U900 ( .A0(n103), .A1(n380), .B0(n104), .B1(n383), .C0(n295), .Y(
        in1[2]) );
  NAND2X1 U901 ( .A(read_data1_out[2]), .B(n389), .Y(n295) );
  OAI221XL U902 ( .A0(n136), .A1(n380), .B0(n137), .B1(n388), .C0(n306), .Y(
        in1[1]) );
  NAND2X1 U903 ( .A(read_data1_out[1]), .B(n390), .Y(n306) );
  OAI221XL U904 ( .A0(n136), .A1(n407), .B0(n408), .B1(n137), .C0(n138), .Y(
        source2[1]) );
  AOI22X1 U905 ( .A0(read_data2_out[1]), .A1(n353), .B0(ext_reg_out[1]), .B1(
        sel_in2_out), .Y(n138) );
  OAI2BB1X1 U906 ( .A0N(next_pc[0]), .A1N(stall), .B0(n351), .Y(N35) );
  AOI22X1 U907 ( .A0(N92), .A1(n361), .B0(pc_shift[0]), .B1(n372), .Y(n351) );
  OAI221XL U908 ( .A0(n169), .A1(n380), .B0(n170), .B1(n383), .C0(n317), .Y(
        in1[0]) );
  NAND2X1 U909 ( .A(read_data1_out[0]), .B(n389), .Y(n317) );
  OAI221XL U910 ( .A0(n88), .A1(n406), .B0(n408), .B1(n89), .C0(n90), .Y(
        source2[5]) );
  AOI22X1 U911 ( .A0(read_data2_out[5]), .A1(n353), .B0(ext_reg_out[5]), .B1(
        sel_in2_out), .Y(n90) );
  OAI2BB1X1 U912 ( .A0N(next_pc[1]), .A1N(stall), .B0(n350), .Y(N36) );
  AOI22X1 U913 ( .A0(N93), .A1(n361), .B0(pc_shift[1]), .B1(n373), .Y(n350) );
  OAI2BB1X1 U914 ( .A0N(next_pc[2]), .A1N(stall), .B0(n349), .Y(N37) );
  AOI22X1 U915 ( .A0(N94), .A1(n361), .B0(pc_shift[2]), .B1(n373), .Y(n349) );
  OAI2BB1X1 U916 ( .A0N(next_pc[3]), .A1N(stall), .B0(n348), .Y(N38) );
  AOI22X1 U917 ( .A0(N95), .A1(n361), .B0(pc_shift[3]), .B1(n374), .Y(n348) );
  OAI2BB1X1 U918 ( .A0N(next_pc[4]), .A1N(stall), .B0(n347), .Y(N39) );
  AOI22X1 U919 ( .A0(N96), .A1(n364), .B0(pc_shift[4]), .B1(n373), .Y(n347) );
  OAI2BB1X1 U920 ( .A0N(next_pc[5]), .A1N(stall), .B0(n346), .Y(N40) );
  AOI22X1 U921 ( .A0(N97), .A1(n367), .B0(pc_shift[5]), .B1(n374), .Y(n346) );
  OAI2BB1X1 U922 ( .A0N(next_pc[6]), .A1N(stall), .B0(n345), .Y(N41) );
  AOI22X1 U923 ( .A0(N98), .A1(n363), .B0(pc_shift[6]), .B1(n376), .Y(n345) );
  OAI2BB1X1 U924 ( .A0N(next_pc[7]), .A1N(stall), .B0(n344), .Y(N42) );
  AOI22X1 U925 ( .A0(N99), .A1(n363), .B0(pc_shift[7]), .B1(n374), .Y(n344) );
  OAI2BB1X1 U926 ( .A0N(next_pc[8]), .A1N(stall), .B0(n343), .Y(N43) );
  AOI22X1 U927 ( .A0(N100), .A1(n364), .B0(pc_shift[8]), .B1(n376), .Y(n343)
         );
  OAI2BB1X1 U928 ( .A0N(next_pc[9]), .A1N(stall), .B0(n342), .Y(N44) );
  AOI22X1 U929 ( .A0(N101), .A1(n364), .B0(pc_shift[9]), .B1(n378), .Y(n342)
         );
  OAI2BB1X1 U930 ( .A0N(next_pc[10]), .A1N(stall), .B0(n341), .Y(N45) );
  AOI22X1 U931 ( .A0(N102), .A1(n364), .B0(pc_shift[10]), .B1(n376), .Y(n341)
         );
  OAI2BB1X1 U932 ( .A0N(next_pc[11]), .A1N(stall), .B0(n340), .Y(N46) );
  AOI22X1 U933 ( .A0(N103), .A1(n365), .B0(pc_shift[11]), .B1(n379), .Y(n340)
         );
  OAI2BB1X1 U934 ( .A0N(next_pc[14]), .A1N(stall), .B0(n337), .Y(N49) );
  AOI22X1 U935 ( .A0(N106), .A1(n364), .B0(pc_shift[14]), .B1(n376), .Y(n337)
         );
  OAI2BB1X1 U936 ( .A0N(next_pc[15]), .A1N(stall), .B0(n336), .Y(N50) );
  AOI22X1 U937 ( .A0(N107), .A1(n365), .B0(pc_shift[15]), .B1(n320), .Y(n336)
         );
  OAI2BB1X1 U938 ( .A0N(next_pc[22]), .A1N(stall), .B0(n329), .Y(N57) );
  AOI22X1 U939 ( .A0(N114), .A1(n361), .B0(pc_shift[22]), .B1(n372), .Y(n329)
         );
  OAI2BB1X1 U940 ( .A0N(next_pc[23]), .A1N(stall), .B0(n328), .Y(N58) );
  AOI22X1 U941 ( .A0(N115), .A1(n358), .B0(pc_shift[23]), .B1(n373), .Y(n328)
         );
  OAI2BB1X1 U942 ( .A0N(next_pc[24]), .A1N(stall), .B0(n327), .Y(N59) );
  AOI22X1 U943 ( .A0(N116), .A1(n363), .B0(pc_shift[24]), .B1(n372), .Y(n327)
         );
  OAI2BB1X1 U944 ( .A0N(next_pc[25]), .A1N(stall), .B0(n326), .Y(N60) );
  AOI22X1 U945 ( .A0(N117), .A1(n358), .B0(pc_shift[25]), .B1(n374), .Y(n326)
         );
  OAI2BB1X1 U946 ( .A0N(next_pc[26]), .A1N(stall), .B0(n325), .Y(N61) );
  AOI22X1 U947 ( .A0(N118), .A1(n368), .B0(pc_shift[26]), .B1(n374), .Y(n325)
         );
  OAI2BB1X1 U948 ( .A0N(next_pc[27]), .A1N(stall), .B0(n324), .Y(N62) );
  AOI22X1 U949 ( .A0(N119), .A1(n319), .B0(pc_shift[27]), .B1(n372), .Y(n324)
         );
  OAI2BB1X1 U950 ( .A0N(next_pc[28]), .A1N(stall), .B0(n323), .Y(N63) );
  AOI22X1 U951 ( .A0(N120), .A1(n363), .B0(pc_shift[28]), .B1(n372), .Y(n323)
         );
  OAI2BB1X1 U952 ( .A0N(next_pc[29]), .A1N(stall), .B0(n322), .Y(N64) );
  AOI22X1 U953 ( .A0(N121), .A1(n363), .B0(pc_shift[29]), .B1(n370), .Y(n322)
         );
  OAI2BB1X1 U954 ( .A0N(next_pc[30]), .A1N(stall), .B0(n321), .Y(N65) );
  AOI22X1 U955 ( .A0(N122), .A1(n365), .B0(pc_shift[30]), .B1(n373), .Y(n321)
         );
  OAI2BB1X1 U956 ( .A0N(stall), .A1N(next_pc[31]), .B0(n318), .Y(N66) );
  AOI22X1 U957 ( .A0(N123), .A1(n365), .B0(pc_shift[31]), .B1(n376), .Y(n318)
         );
  OAI2BB1X1 U958 ( .A0N(next_pc[12]), .A1N(stall), .B0(n339), .Y(N47) );
  AOI22X1 U959 ( .A0(N104), .A1(n367), .B0(pc_shift[12]), .B1(n378), .Y(n339)
         );
  OAI2BB1X1 U960 ( .A0N(next_pc[13]), .A1N(stall), .B0(n338), .Y(N48) );
  AOI22X1 U961 ( .A0(N105), .A1(n367), .B0(pc_shift[13]), .B1(n378), .Y(n338)
         );
  OAI2BB1X1 U962 ( .A0N(next_pc[16]), .A1N(stall), .B0(n335), .Y(N51) );
  AOI22X1 U963 ( .A0(N108), .A1(n367), .B0(pc_shift[16]), .B1(n378), .Y(n335)
         );
  OAI2BB1X1 U964 ( .A0N(next_pc[17]), .A1N(stall), .B0(n334), .Y(N52) );
  AOI22X1 U965 ( .A0(N109), .A1(n368), .B0(pc_shift[17]), .B1(n378), .Y(n334)
         );
  OAI221XL U966 ( .A0(n169), .A1(n403), .B0(n408), .B1(n170), .C0(n171), .Y(
        source2[0]) );
  AOI22X1 U967 ( .A0(read_data2_out[0]), .A1(n353), .B0(ext_reg_out[0]), .B1(
        sel_in2_out), .Y(n171) );
  INVX1 U968 ( .A(sel_in2_out), .Y(n424) );
  INVX1 U969 ( .A(sel_wb_reg2_out), .Y(n412) );
  INVX1 U970 ( .A(sel_wb_reg2_out), .Y(n413) );
  OAI221XL U971 ( .A0(n109), .A1(n404), .B0(n408), .B1(n110), .C0(n111), .Y(
        source2[28]) );
  AOI22X1 U972 ( .A0(read_data2_out[28]), .A1(n353), .B0(ext_reg_out[28]), 
        .B1(sel_in2_out), .Y(n111) );
  OAI221XL U973 ( .A0(n112), .A1(n404), .B0(n408), .B1(n113), .C0(n114), .Y(
        source2[27]) );
  AOI22X1 U974 ( .A0(read_data2_out[27]), .A1(n353), .B0(ext_reg_out[27]), 
        .B1(sel_in2_out), .Y(n114) );
  OAI221XL U975 ( .A0(n115), .A1(n404), .B0(n408), .B1(n116), .C0(n117), .Y(
        source2[26]) );
  AOI22X1 U976 ( .A0(read_data2_out[26]), .A1(n353), .B0(ext_reg_out[26]), 
        .B1(sel_in2_out), .Y(n117) );
  OAI221XL U977 ( .A0(n127), .A1(n404), .B0(n408), .B1(n128), .C0(n129), .Y(
        source2[22]) );
  AOI22X1 U978 ( .A0(read_data2_out[22]), .A1(n353), .B0(ext_reg_out[22]), 
        .B1(sel_in2_out), .Y(n129) );
  OAI221XL U979 ( .A0(n118), .A1(n404), .B0(n408), .B1(n119), .C0(n120), .Y(
        source2[25]) );
  AOI22X1 U980 ( .A0(read_data2_out[25]), .A1(n353), .B0(ext_reg_out[25]), 
        .B1(sel_in2_out), .Y(n120) );
  OAI221XL U981 ( .A0(n106), .A1(n404), .B0(n408), .B1(n107), .C0(n108), .Y(
        source2[29]) );
  AOI22X1 U982 ( .A0(read_data2_out[29]), .A1(n353), .B0(ext_reg_out[29]), 
        .B1(sel_in2_out), .Y(n108) );
  OAI221XL U983 ( .A0(n100), .A1(n404), .B0(n408), .B1(n101), .C0(n102), .Y(
        source2[30]) );
  AOI22X1 U984 ( .A0(read_data2_out[30]), .A1(n353), .B0(ext_reg_out[30]), 
        .B1(sel_in2_out), .Y(n102) );
  OAI221XL U985 ( .A0(n121), .A1(n404), .B0(n408), .B1(n122), .C0(n123), .Y(
        source2[24]) );
  AOI22X1 U986 ( .A0(read_data2_out[24]), .A1(n353), .B0(ext_reg_out[24]), 
        .B1(sel_in2_out), .Y(n123) );
  OAI221XL U987 ( .A0(n142), .A1(n404), .B0(n408), .B1(n143), .C0(n144), .Y(
        source2[18]) );
  AOI22X1 U988 ( .A0(read_data2_out[18]), .A1(n353), .B0(ext_reg_out[18]), 
        .B1(sel_in2_out), .Y(n144) );
  OAI221XL U989 ( .A0(n148), .A1(n405), .B0(n408), .B1(n149), .C0(n150), .Y(
        source2[16]) );
  AOI22X1 U990 ( .A0(read_data2_out[16]), .A1(n353), .B0(ext_reg_out[16]), 
        .B1(sel_in2_out), .Y(n150) );
  OAI221XL U991 ( .A0(n130), .A1(n404), .B0(n408), .B1(n131), .C0(n132), .Y(
        source2[21]) );
  AOI22X1 U992 ( .A0(read_data2_out[21]), .A1(n353), .B0(ext_reg_out[21]), 
        .B1(sel_in2_out), .Y(n132) );
  OAI221XL U993 ( .A0(n160), .A1(n404), .B0(n408), .B1(n161), .C0(n162), .Y(
        source2[12]) );
  AOI22X1 U994 ( .A0(read_data2_out[12]), .A1(n353), .B0(ext_reg_out[12]), 
        .B1(sel_in2_out), .Y(n162) );
  OAI221XL U995 ( .A0(n139), .A1(n404), .B0(n408), .B1(n140), .C0(n141), .Y(
        source2[19]) );
  AOI22X1 U996 ( .A0(read_data2_out[19]), .A1(n353), .B0(ext_reg_out[19]), 
        .B1(sel_in2_out), .Y(n141) );
  OAI221XL U997 ( .A0(n133), .A1(n404), .B0(n408), .B1(n134), .C0(n135), .Y(
        source2[20]) );
  AOI22X1 U998 ( .A0(read_data2_out[20]), .A1(n353), .B0(ext_reg_out[20]), 
        .B1(sel_in2_out), .Y(n135) );
  OAI221XL U999 ( .A0(n145), .A1(n406), .B0(n408), .B1(n146), .C0(n147), .Y(
        source2[17]) );
  AOI22X1 U1000 ( .A0(read_data2_out[17]), .A1(n353), .B0(ext_reg_out[17]), 
        .B1(sel_in2_out), .Y(n147) );
  OAI221XL U1001 ( .A0(n151), .A1(n404), .B0(n408), .B1(n152), .C0(n153), .Y(
        source2[15]) );
  AOI22X1 U1002 ( .A0(read_data2_out[15]), .A1(n353), .B0(ext_reg_out[15]), 
        .B1(sel_in2_out), .Y(n153) );
  OAI221XL U1003 ( .A0(n154), .A1(n380), .B0(n155), .B1(n386), .C0(n312), .Y(
        in1[14]) );
  NAND2X1 U1004 ( .A(read_data1_out[14]), .B(n390), .Y(n312) );
  OAI221XL U1005 ( .A0(n137), .A1(n391), .B0(n256), .B1(n392), .C0(n257), .Y(
        read_data1_in[1]) );
  AOI22X1 U1006 ( .A0(n394), .A1(write_data[1]), .B0(read_data1[1]), .B1(n396), 
        .Y(n257) );
  AOI22X1 U1007 ( .A0(n416), .A1(alu_result_reg_out[9]), .B0(data_out_out[9]), 
        .B1(n420), .Y(n73) );
  AOI22X1 U1008 ( .A0(alu_result_reg_out[10]), .A1(n414), .B0(data_out_out[10]), .B1(n422), .Y(n166) );
  AOI22X1 U1009 ( .A0(alu_result_reg_out[11]), .A1(n414), .B0(data_out_out[11]), .B1(n420), .Y(n163) );
  AOI22X1 U1010 ( .A0(alu_result_reg_out[12]), .A1(n414), .B0(data_out_out[12]), .B1(n420), .Y(n160) );
  AOI22X1 U1011 ( .A0(alu_result_reg_out[13]), .A1(n414), .B0(data_out_out[13]), .B1(n420), .Y(n157) );
  AOI22X1 U1012 ( .A0(alu_result_reg_out[14]), .A1(n414), .B0(data_out_out[14]), .B1(n420), .Y(n154) );
  AOI22X1 U1013 ( .A0(alu_result_reg_out[15]), .A1(n414), .B0(data_out_out[15]), .B1(n420), .Y(n151) );
  AOI22X1 U1014 ( .A0(alu_result_reg_out[16]), .A1(n414), .B0(data_out_out[16]), .B1(n420), .Y(n148) );
  AOI22X1 U1015 ( .A0(alu_result_reg_out[17]), .A1(n414), .B0(data_out_out[17]), .B1(n420), .Y(n145) );
  AOI22X1 U1016 ( .A0(alu_result_reg_out[18]), .A1(n414), .B0(data_out_out[18]), .B1(n420), .Y(n142) );
  AOI22X1 U1017 ( .A0(alu_result_reg_out[19]), .A1(n414), .B0(data_out_out[19]), .B1(n421), .Y(n139) );
  AOI22X1 U1018 ( .A0(alu_result_reg_out[20]), .A1(n415), .B0(data_out_out[20]), .B1(n420), .Y(n133) );
  AOI22X1 U1019 ( .A0(alu_result_reg_out[21]), .A1(n415), .B0(data_out_out[21]), .B1(n420), .Y(n130) );
  AOI22X1 U1020 ( .A0(alu_result_reg_out[22]), .A1(n415), .B0(data_out_out[22]), .B1(n420), .Y(n127) );
  AOI22X1 U1021 ( .A0(alu_result_reg_out[23]), .A1(n415), .B0(data_out_out[23]), .B1(n420), .Y(n124) );
  AOI22X1 U1022 ( .A0(alu_result_reg_out[24]), .A1(n415), .B0(data_out_out[24]), .B1(n420), .Y(n121) );
  AOI22X1 U1023 ( .A0(alu_result_reg_out[25]), .A1(n415), .B0(data_out_out[25]), .B1(n420), .Y(n118) );
  AOI22X1 U1024 ( .A0(alu_result_reg_out[26]), .A1(n415), .B0(data_out_out[26]), .B1(n420), .Y(n115) );
  AOI22X1 U1025 ( .A0(alu_result_reg_out[27]), .A1(n415), .B0(data_out_out[27]), .B1(n420), .Y(n112) );
  AOI22X1 U1026 ( .A0(alu_result_reg_out[28]), .A1(n415), .B0(data_out_out[28]), .B1(n420), .Y(n109) );
  AOI22X1 U1027 ( .A0(alu_result_reg_out[29]), .A1(n415), .B0(data_out_out[29]), .B1(n420), .Y(n106) );
  AOI22X1 U1028 ( .A0(alu_result_reg_out[30]), .A1(n415), .B0(data_out_out[30]), .B1(n419), .Y(n100) );
  OAI221XL U1029 ( .A0(n169), .A1(n356), .B0(n170), .B1(n357), .C0(n209), .Y(
        read_data3_in[0]) );
  AOI22X1 U1030 ( .A0(result[0]), .A1(n354), .B0(read_data3[0]), .B1(n355), 
        .Y(n209) );
  OAI221XL U1031 ( .A0(n170), .A1(n391), .B0(n278), .B1(n392), .C0(n279), .Y(
        read_data1_in[0]) );
  AOI22X1 U1032 ( .A0(n394), .A1(write_data[0]), .B0(read_data1[0]), .B1(n395), 
        .Y(n279) );
  OAI221XL U1033 ( .A0(n103), .A1(n356), .B0(n104), .B1(n357), .C0(n187), .Y(
        read_data3_in[2]) );
  AOI22X1 U1034 ( .A0(result[2]), .A1(n354), .B0(read_data3[2]), .B1(n355), 
        .Y(n187) );
  OAI221XL U1035 ( .A0(n94), .A1(n356), .B0(n95), .B1(n357), .C0(n184), .Y(
        read_data3_in[3]) );
  AOI22X1 U1036 ( .A0(result[3]), .A1(n354), .B0(read_data3[3]), .B1(n355), 
        .Y(n184) );
  OAI221XL U1037 ( .A0(n91), .A1(n356), .B0(n92), .B1(n357), .C0(n183), .Y(
        read_data3_in[4]) );
  AOI22X1 U1038 ( .A0(result[4]), .A1(n354), .B0(read_data3[4]), .B1(n355), 
        .Y(n183) );
  OAI221XL U1039 ( .A0(n88), .A1(n356), .B0(n89), .B1(n357), .C0(n182), .Y(
        read_data3_in[5]) );
  AOI22X1 U1040 ( .A0(result[5]), .A1(n354), .B0(read_data3[5]), .B1(n355), 
        .Y(n182) );
  OAI221XL U1041 ( .A0(n85), .A1(n356), .B0(n86), .B1(n357), .C0(n181), .Y(
        read_data3_in[6]) );
  AOI22X1 U1042 ( .A0(result[6]), .A1(n354), .B0(read_data3[6]), .B1(n355), 
        .Y(n181) );
  OAI221XL U1043 ( .A0(n82), .A1(n356), .B0(n83), .B1(n357), .C0(n180), .Y(
        read_data3_in[7]) );
  AOI22X1 U1044 ( .A0(result[7]), .A1(n354), .B0(read_data3[7]), .B1(n355), 
        .Y(n180) );
  OAI221XL U1045 ( .A0(n79), .A1(n356), .B0(n80), .B1(n357), .C0(n179), .Y(
        read_data3_in[8]) );
  AOI22X1 U1046 ( .A0(result[8]), .A1(n354), .B0(read_data3[8]), .B1(n355), 
        .Y(n179) );
  OAI221XL U1047 ( .A0(n73), .A1(n356), .B0(n76), .B1(n357), .C0(n176), .Y(
        read_data3_in[9]) );
  AOI22X1 U1048 ( .A0(result[9]), .A1(n354), .B0(read_data3[9]), .B1(n355), 
        .Y(n176) );
  OAI221XL U1049 ( .A0(n166), .A1(n356), .B0(n167), .B1(n357), .C0(n208), .Y(
        read_data3_in[10]) );
  AOI22X1 U1050 ( .A0(result[10]), .A1(n354), .B0(read_data3[10]), .B1(n355), 
        .Y(n208) );
  OAI221XL U1051 ( .A0(n163), .A1(n356), .B0(n164), .B1(n357), .C0(n207), .Y(
        read_data3_in[11]) );
  AOI22X1 U1052 ( .A0(result[11]), .A1(n354), .B0(read_data3[11]), .B1(n355), 
        .Y(n207) );
  OAI221XL U1053 ( .A0(n160), .A1(n356), .B0(n161), .B1(n357), .C0(n206), .Y(
        read_data3_in[12]) );
  AOI22X1 U1054 ( .A0(result[12]), .A1(n354), .B0(read_data3[12]), .B1(n355), 
        .Y(n206) );
  OAI221XL U1055 ( .A0(n157), .A1(n356), .B0(n158), .B1(n357), .C0(n205), .Y(
        read_data3_in[13]) );
  AOI22X1 U1056 ( .A0(result[13]), .A1(n354), .B0(read_data3[13]), .B1(n355), 
        .Y(n205) );
  OAI221XL U1057 ( .A0(n154), .A1(n356), .B0(n155), .B1(n357), .C0(n204), .Y(
        read_data3_in[14]) );
  AOI22X1 U1058 ( .A0(result[14]), .A1(n354), .B0(read_data3[14]), .B1(n355), 
        .Y(n204) );
  OAI221XL U1059 ( .A0(n151), .A1(n356), .B0(n152), .B1(n357), .C0(n203), .Y(
        read_data3_in[15]) );
  AOI22X1 U1060 ( .A0(result[15]), .A1(n354), .B0(read_data3[15]), .B1(n355), 
        .Y(n203) );
  OAI221XL U1061 ( .A0(n148), .A1(n356), .B0(n149), .B1(n357), .C0(n202), .Y(
        read_data3_in[16]) );
  AOI22X1 U1062 ( .A0(result[16]), .A1(n354), .B0(read_data3[16]), .B1(n355), 
        .Y(n202) );
  OAI221XL U1063 ( .A0(n145), .A1(n356), .B0(n146), .B1(n357), .C0(n201), .Y(
        read_data3_in[17]) );
  AOI22X1 U1064 ( .A0(result[17]), .A1(n354), .B0(read_data3[17]), .B1(n355), 
        .Y(n201) );
  OAI221XL U1065 ( .A0(n142), .A1(n356), .B0(n143), .B1(n357), .C0(n200), .Y(
        read_data3_in[18]) );
  AOI22X1 U1066 ( .A0(result[18]), .A1(n354), .B0(read_data3[18]), .B1(n355), 
        .Y(n200) );
  OAI221XL U1067 ( .A0(n139), .A1(n356), .B0(n140), .B1(n357), .C0(n199), .Y(
        read_data3_in[19]) );
  AOI22X1 U1068 ( .A0(result[19]), .A1(n354), .B0(read_data3[19]), .B1(n355), 
        .Y(n199) );
  OAI221XL U1069 ( .A0(n133), .A1(n356), .B0(n134), .B1(n357), .C0(n197), .Y(
        read_data3_in[20]) );
  AOI22X1 U1070 ( .A0(result[20]), .A1(n354), .B0(read_data3[20]), .B1(n355), 
        .Y(n197) );
  OAI221XL U1071 ( .A0(n104), .A1(n391), .B0(n234), .B1(n392), .C0(n235), .Y(
        read_data1_in[2]) );
  AOI22X1 U1072 ( .A0(n393), .A1(write_data[2]), .B0(read_data1[2]), .B1(n395), 
        .Y(n235) );
  OAI221XL U1073 ( .A0(n95), .A1(n391), .B0(n228), .B1(n392), .C0(n229), .Y(
        read_data1_in[3]) );
  AOI22X1 U1074 ( .A0(n393), .A1(write_data[3]), .B0(read_data1[3]), .B1(n395), 
        .Y(n229) );
  OAI221XL U1075 ( .A0(n92), .A1(n391), .B0(n226), .B1(n392), .C0(n227), .Y(
        read_data1_in[4]) );
  AOI22X1 U1076 ( .A0(n393), .A1(write_data[4]), .B0(read_data1[4]), .B1(n395), 
        .Y(n227) );
  OAI221XL U1077 ( .A0(n89), .A1(n391), .B0(n224), .B1(n392), .C0(n225), .Y(
        read_data1_in[5]) );
  AOI22X1 U1078 ( .A0(n393), .A1(write_data[5]), .B0(read_data1[5]), .B1(n395), 
        .Y(n225) );
  OAI221XL U1079 ( .A0(n86), .A1(n391), .B0(n222), .B1(n392), .C0(n223), .Y(
        read_data1_in[6]) );
  AOI22X1 U1080 ( .A0(n393), .A1(write_data[6]), .B0(read_data1[6]), .B1(n396), 
        .Y(n223) );
  OAI221XL U1081 ( .A0(n83), .A1(n391), .B0(n220), .B1(n392), .C0(n221), .Y(
        read_data1_in[7]) );
  AOI22X1 U1082 ( .A0(n393), .A1(write_data[7]), .B0(read_data1[7]), .B1(n396), 
        .Y(n221) );
  OAI221XL U1083 ( .A0(n80), .A1(n391), .B0(n218), .B1(n392), .C0(n219), .Y(
        read_data1_in[8]) );
  AOI22X1 U1084 ( .A0(n393), .A1(write_data[8]), .B0(read_data1[8]), .B1(n396), 
        .Y(n219) );
  OAI221XL U1085 ( .A0(n76), .A1(n391), .B0(n213), .B1(n392), .C0(n215), .Y(
        read_data1_in[9]) );
  AOI22X1 U1086 ( .A0(n394), .A1(write_data[9]), .B0(read_data1[9]), .B1(n396), 
        .Y(n215) );
  OAI221XL U1087 ( .A0(n167), .A1(n391), .B0(n276), .B1(n392), .C0(n277), .Y(
        read_data1_in[10]) );
  AOI22X1 U1088 ( .A0(n394), .A1(write_data[10]), .B0(read_data1[10]), .B1(
        n395), .Y(n277) );
  OAI221XL U1089 ( .A0(n164), .A1(n391), .B0(n274), .B1(n392), .C0(n275), .Y(
        read_data1_in[11]) );
  AOI22X1 U1090 ( .A0(n394), .A1(write_data[11]), .B0(read_data1[11]), .B1(
        n395), .Y(n275) );
  OAI221XL U1091 ( .A0(n161), .A1(n391), .B0(n272), .B1(n392), .C0(n273), .Y(
        read_data1_in[12]) );
  AOI22X1 U1092 ( .A0(n394), .A1(write_data[12]), .B0(read_data1[12]), .B1(
        n395), .Y(n273) );
  OAI221XL U1093 ( .A0(n158), .A1(n391), .B0(n270), .B1(n392), .C0(n271), .Y(
        read_data1_in[13]) );
  AOI22X1 U1094 ( .A0(n394), .A1(write_data[13]), .B0(read_data1[13]), .B1(
        n395), .Y(n271) );
  OAI221XL U1095 ( .A0(n155), .A1(n391), .B0(n268), .B1(n392), .C0(n269), .Y(
        read_data1_in[14]) );
  AOI22X1 U1096 ( .A0(n394), .A1(write_data[14]), .B0(read_data1[14]), .B1(
        n395), .Y(n269) );
  OAI221XL U1097 ( .A0(n152), .A1(n391), .B0(n266), .B1(n392), .C0(n267), .Y(
        read_data1_in[15]) );
  AOI22X1 U1098 ( .A0(n394), .A1(write_data[15]), .B0(read_data1[15]), .B1(
        n396), .Y(n267) );
  OAI221XL U1099 ( .A0(n149), .A1(n391), .B0(n264), .B1(n392), .C0(n265), .Y(
        read_data1_in[16]) );
  AOI22X1 U1100 ( .A0(n394), .A1(write_data[16]), .B0(read_data1[16]), .B1(
        n396), .Y(n265) );
  OAI221XL U1101 ( .A0(n146), .A1(n391), .B0(n262), .B1(n392), .C0(n263), .Y(
        read_data1_in[17]) );
  AOI22X1 U1102 ( .A0(n394), .A1(write_data[17]), .B0(read_data1[17]), .B1(
        n396), .Y(n263) );
  OAI221XL U1103 ( .A0(n143), .A1(n391), .B0(n260), .B1(n392), .C0(n261), .Y(
        read_data1_in[18]) );
  AOI22X1 U1104 ( .A0(n394), .A1(write_data[18]), .B0(read_data1[18]), .B1(
        n396), .Y(n261) );
  OAI221XL U1105 ( .A0(n140), .A1(n391), .B0(n258), .B1(n392), .C0(n259), .Y(
        read_data1_in[19]) );
  AOI22X1 U1106 ( .A0(n394), .A1(write_data[19]), .B0(read_data1[19]), .B1(
        n396), .Y(n259) );
  OAI221XL U1107 ( .A0(n134), .A1(n391), .B0(n254), .B1(n392), .C0(n255), .Y(
        read_data1_in[20]) );
  AOI22X1 U1108 ( .A0(n394), .A1(write_data[20]), .B0(read_data1[20]), .B1(
        n217), .Y(n255) );
  OAI221XL U1109 ( .A0(n136), .A1(n356), .B0(n137), .B1(n357), .C0(n198), .Y(
        read_data3_in[1]) );
  AOI22X1 U1110 ( .A0(result[1]), .A1(n354), .B0(read_data3[1]), .B1(n355), 
        .Y(n198) );
  OAI2BB2X1 U1111 ( .B0(sel_alu_out), .B1(n246), .A0N(ext_reg_out[24]), .A1N(
        sel_alu_out), .Y(alu_result[24]) );
  OAI2BB2X1 U1112 ( .B0(sel_alu_out), .B1(n244), .A0N(ext_reg_out[25]), .A1N(
        sel_alu_out), .Y(alu_result[25]) );
  OAI2BB2X1 U1113 ( .B0(sel_alu_out), .B1(n242), .A0N(ext_reg_out[26]), .A1N(
        sel_alu_out), .Y(alu_result[26]) );
  OAI2BB2X1 U1114 ( .B0(sel_alu_out), .B1(n240), .A0N(ext_reg_out[27]), .A1N(
        sel_alu_out), .Y(alu_result[27]) );
  OAI2BB2X1 U1115 ( .B0(sel_alu_out), .B1(n238), .A0N(ext_reg_out[28]), .A1N(
        sel_alu_out), .Y(alu_result[28]) );
  OAI2BB2X1 U1116 ( .B0(sel_alu_out), .B1(n236), .A0N(ext_reg_out[29]), .A1N(
        sel_alu_out), .Y(alu_result[29]) );
  OAI2BB2X1 U1117 ( .B0(sel_alu_out), .B1(n232), .A0N(ext_reg_out[30]), .A1N(
        sel_alu_out), .Y(alu_result[30]) );
  OAI2BB2X1 U1118 ( .B0(sel_alu_out), .B1(n230), .A0N(ext_reg_out[31]), .A1N(
        sel_alu_out), .Y(alu_result[31]) );
  OAI221XL U1119 ( .A0(n163), .A1(n404), .B0(n408), .B1(n164), .C0(n165), .Y(
        source2[11]) );
  AOI22X1 U1120 ( .A0(read_data2_out[11]), .A1(n353), .B0(ext_reg_out[11]), 
        .B1(sel_in2_out), .Y(n165) );
  OAI221XL U1121 ( .A0(n157), .A1(n404), .B0(n408), .B1(n158), .C0(n159), .Y(
        source2[13]) );
  AOI22X1 U1122 ( .A0(read_data2_out[13]), .A1(n353), .B0(ext_reg_out[13]), 
        .B1(sel_in2_out), .Y(n159) );
  OAI221XL U1123 ( .A0(n154), .A1(n404), .B0(n408), .B1(n155), .C0(n156), .Y(
        source2[14]) );
  AOI22X1 U1124 ( .A0(read_data2_out[14]), .A1(n353), .B0(ext_reg_out[14]), 
        .B1(sel_in2_out), .Y(n156) );
  OAI221XL U1125 ( .A0(n124), .A1(n407), .B0(n408), .B1(n125), .C0(n126), .Y(
        source2[23]) );
  AOI22X1 U1126 ( .A0(read_data2_out[23]), .A1(n353), .B0(ext_reg_out[23]), 
        .B1(sel_in2_out), .Y(n126) );
  OAI221XL U1127 ( .A0(n97), .A1(n404), .B0(n408), .B1(n98), .C0(n99), .Y(
        source2[31]) );
  AOI22X1 U1128 ( .A0(read_data2_out[31]), .A1(n353), .B0(ext_reg_out[31]), 
        .B1(sel_in2_out), .Y(n99) );
  INVX1 U1129 ( .A(alu_result_out[3]), .Y(n95) );
  INVX1 U1130 ( .A(alu_result_out[4]), .Y(n92) );
  INVX1 U1131 ( .A(alu_result_out[5]), .Y(n89) );
  INVX1 U1132 ( .A(alu_result_out[6]), .Y(n86) );
  INVX1 U1133 ( .A(alu_result_out[7]), .Y(n83) );
  INVX1 U1134 ( .A(alu_result_out[8]), .Y(n80) );
  INVX1 U1135 ( .A(alu_result_out[9]), .Y(n76) );
  INVX1 U1136 ( .A(alu_result_out[10]), .Y(n167) );
  INVX1 U1137 ( .A(alu_result_out[11]), .Y(n164) );
  INVX1 U1138 ( .A(alu_result_out[12]), .Y(n161) );
  INVX1 U1139 ( .A(alu_result_out[13]), .Y(n158) );
  INVX1 U1140 ( .A(alu_result_out[14]), .Y(n155) );
  OAI221XL U1141 ( .A0(n151), .A1(n380), .B0(n152), .B1(n387), .C0(n311), .Y(
        in1[15]) );
  NAND2X1 U1142 ( .A(read_data1_out[15]), .B(n389), .Y(n311) );
  OAI221XL U1143 ( .A0(n148), .A1(n380), .B0(n149), .B1(n387), .C0(n310), .Y(
        in1[16]) );
  NAND2X1 U1144 ( .A(read_data1_out[16]), .B(n390), .Y(n310) );
  OAI221XL U1145 ( .A0(n166), .A1(n380), .B0(n167), .B1(n387), .C0(n316), .Y(
        in1[10]) );
  NAND2X1 U1146 ( .A(read_data1_out[10]), .B(n390), .Y(n316) );
  OAI221XL U1147 ( .A0(n163), .A1(n380), .B0(n164), .B1(n387), .C0(n315), .Y(
        in1[11]) );
  NAND2X1 U1148 ( .A(read_data1_out[11]), .B(n389), .Y(n315) );
  OAI221XL U1149 ( .A0(n160), .A1(n380), .B0(n161), .B1(n384), .C0(n314), .Y(
        in1[12]) );
  NAND2X1 U1150 ( .A(read_data1_out[12]), .B(n390), .Y(n314) );
  OAI221XL U1151 ( .A0(n157), .A1(n380), .B0(n158), .B1(n385), .C0(n313), .Y(
        in1[13]) );
  NAND2X1 U1152 ( .A(read_data1_out[13]), .B(n389), .Y(n313) );
  OAI221XL U1153 ( .A0(n145), .A1(n380), .B0(n146), .B1(n387), .C0(n309), .Y(
        in1[17]) );
  NAND2X1 U1154 ( .A(read_data1_out[17]), .B(n389), .Y(n309) );
  OAI221XL U1155 ( .A0(n142), .A1(n380), .B0(n143), .B1(n387), .C0(n308), .Y(
        in1[18]) );
  NAND2X1 U1156 ( .A(read_data1_out[18]), .B(n390), .Y(n308) );
  OAI221XL U1157 ( .A0(n139), .A1(n380), .B0(n140), .B1(n387), .C0(n307), .Y(
        in1[19]) );
  NAND2X1 U1158 ( .A(read_data1_out[19]), .B(n389), .Y(n307) );
  OAI221XL U1159 ( .A0(n133), .A1(n380), .B0(n134), .B1(n387), .C0(n305), .Y(
        in1[20]) );
  NAND2X1 U1160 ( .A(read_data1_out[20]), .B(n389), .Y(n305) );
  OAI221XL U1161 ( .A0(n106), .A1(n380), .B0(n107), .B1(n386), .C0(n296), .Y(
        in1[29]) );
  NAND2X1 U1162 ( .A(read_data1_out[29]), .B(n390), .Y(n296) );
  AOI22X1 U1163 ( .A0(alu_result_reg_out[31]), .A1(n416), .B0(data_out_out[31]), .B1(n418), .Y(n97) );
  OAI2BB2X1 U1164 ( .B0(sel_alu_out), .B1(n222), .A0N(ext_reg_out[6]), .A1N(
        sel_alu_out), .Y(alu_result[6]) );
  OAI2BB2X1 U1165 ( .B0(sel_alu_out), .B1(n220), .A0N(ext_reg_out[7]), .A1N(
        sel_alu_out), .Y(alu_result[7]) );
  OAI2BB2X1 U1166 ( .B0(sel_alu_out), .B1(n218), .A0N(ext_reg_out[8]), .A1N(
        sel_alu_out), .Y(alu_result[8]) );
  OAI2BB2X1 U1167 ( .B0(sel_alu_out), .B1(n213), .A0N(ext_reg_out[9]), .A1N(
        sel_alu_out), .Y(alu_result[9]) );
  OAI2BB2X1 U1168 ( .B0(sel_alu_out), .B1(n276), .A0N(ext_reg_out[10]), .A1N(
        sel_alu_out), .Y(alu_result[10]) );
  OAI2BB2X1 U1169 ( .B0(sel_alu_out), .B1(n274), .A0N(ext_reg_out[11]), .A1N(
        sel_alu_out), .Y(alu_result[11]) );
  OAI2BB2X1 U1170 ( .B0(sel_alu_out), .B1(n272), .A0N(ext_reg_out[12]), .A1N(
        sel_alu_out), .Y(alu_result[12]) );
  OAI2BB2X1 U1171 ( .B0(sel_alu_out), .B1(n270), .A0N(ext_reg_out[13]), .A1N(
        sel_alu_out), .Y(alu_result[13]) );
  OAI2BB2X1 U1172 ( .B0(sel_alu_out), .B1(n268), .A0N(ext_reg_out[14]), .A1N(
        sel_alu_out), .Y(alu_result[14]) );
  OAI2BB2X1 U1173 ( .B0(sel_alu_out), .B1(n266), .A0N(ext_reg_out[15]), .A1N(
        sel_alu_out), .Y(alu_result[15]) );
  OAI2BB2X1 U1174 ( .B0(sel_alu_out), .B1(n264), .A0N(ext_reg_out[16]), .A1N(
        sel_alu_out), .Y(alu_result[16]) );
  OAI2BB2X1 U1175 ( .B0(sel_alu_out), .B1(n262), .A0N(ext_reg_out[17]), .A1N(
        sel_alu_out), .Y(alu_result[17]) );
  OAI2BB2X1 U1176 ( .B0(sel_alu_out), .B1(n260), .A0N(ext_reg_out[18]), .A1N(
        sel_alu_out), .Y(alu_result[18]) );
  OAI2BB2X1 U1177 ( .B0(sel_alu_out), .B1(n258), .A0N(ext_reg_out[19]), .A1N(
        sel_alu_out), .Y(alu_result[19]) );
  OAI2BB2X1 U1178 ( .B0(sel_alu_out), .B1(n254), .A0N(ext_reg_out[20]), .A1N(
        sel_alu_out), .Y(alu_result[20]) );
  OAI2BB2X1 U1179 ( .B0(sel_alu_out), .B1(n252), .A0N(ext_reg_out[21]), .A1N(
        sel_alu_out), .Y(alu_result[21]) );
  OAI2BB2X1 U1180 ( .B0(sel_alu_out), .B1(n250), .A0N(ext_reg_out[22]), .A1N(
        sel_alu_out), .Y(alu_result[22]) );
  OAI2BB2X1 U1181 ( .B0(sel_alu_out), .B1(n248), .A0N(ext_reg_out[23]), .A1N(
        sel_alu_out), .Y(alu_result[23]) );
  OAI2BB2X1 U1182 ( .B0(sel_alu_out), .B1(n278), .A0N(ext_reg_out[0]), .A1N(
        sel_alu_out), .Y(alu_result[0]) );
  OAI2BB2X1 U1183 ( .B0(sel_alu_out), .B1(n256), .A0N(ext_reg_out[1]), .A1N(
        sel_alu_out), .Y(alu_result[1]) );
  OAI2BB2X1 U1184 ( .B0(sel_alu_out), .B1(n234), .A0N(ext_reg_out[2]), .A1N(
        sel_alu_out), .Y(alu_result[2]) );
  OAI2BB2X1 U1185 ( .B0(sel_alu_out), .B1(n228), .A0N(ext_reg_out[3]), .A1N(
        sel_alu_out), .Y(alu_result[3]) );
  OAI2BB2X1 U1186 ( .B0(sel_alu_out), .B1(n226), .A0N(ext_reg_out[4]), .A1N(
        sel_alu_out), .Y(alu_result[4]) );
  OAI2BB2X1 U1187 ( .B0(sel_alu_out), .B1(n224), .A0N(ext_reg_out[5]), .A1N(
        sel_alu_out), .Y(alu_result[5]) );
  OAI221XL U1188 ( .A0(n97), .A1(n380), .B0(n98), .B1(n387), .C0(n293), .Y(
        in1[31]) );
  NAND2X1 U1189 ( .A(read_data1_out[31]), .B(n389), .Y(n293) );
  INVX1 U1190 ( .A(alu_result_out[31]), .Y(n98) );
  INVX1 U1191 ( .A(alu_result_out[15]), .Y(n152) );
  INVX1 U1192 ( .A(alu_result_out[16]), .Y(n149) );
  INVX1 U1193 ( .A(alu_result_out[17]), .Y(n146) );
  INVX1 U1194 ( .A(alu_result_out[18]), .Y(n143) );
  INVX1 U1195 ( .A(alu_result_out[19]), .Y(n140) );
  INVX1 U1196 ( .A(alu_result_out[20]), .Y(n134) );
  INVX1 U1197 ( .A(alu_result_out[21]), .Y(n131) );
  INVX1 U1198 ( .A(alu_result_out[22]), .Y(n128) );
  INVX1 U1199 ( .A(alu_result_out[23]), .Y(n125) );
  INVX1 U1200 ( .A(alu_result_out[24]), .Y(n122) );
  INVX1 U1201 ( .A(alu_result_out[25]), .Y(n119) );
  INVX1 U1202 ( .A(alu_result_out[26]), .Y(n116) );
  INVX1 U1203 ( .A(alu_result_out[27]), .Y(n113) );
  INVX1 U1204 ( .A(alu_result_out[28]), .Y(n110) );
  INVX1 U1205 ( .A(alu_result_out[29]), .Y(n107) );
  INVX1 U1206 ( .A(alu_result_out[30]), .Y(n101) );
  OAI221XL U1207 ( .A0(n100), .A1(n380), .B0(n101), .B1(n387), .C0(n294), .Y(
        in1[30]) );
  NAND2X1 U1208 ( .A(read_data1_out[30]), .B(n390), .Y(n294) );
  OAI221XL U1209 ( .A0(n127), .A1(n380), .B0(n128), .B1(n387), .C0(n303), .Y(
        in1[22]) );
  NAND2X1 U1210 ( .A(read_data1_out[22]), .B(n389), .Y(n303) );
  OAI221XL U1211 ( .A0(n124), .A1(n380), .B0(n125), .B1(n388), .C0(n302), .Y(
        in1[23]) );
  NAND2X1 U1212 ( .A(read_data1_out[23]), .B(n390), .Y(n302) );
  OAI221XL U1213 ( .A0(n121), .A1(n380), .B0(n122), .B1(n387), .C0(n301), .Y(
        in1[24]) );
  NAND2X1 U1214 ( .A(read_data1_out[24]), .B(n389), .Y(n301) );
  OAI221XL U1215 ( .A0(n130), .A1(n380), .B0(n131), .B1(n387), .C0(n304), .Y(
        in1[21]) );
  NAND2X1 U1216 ( .A(read_data1_out[21]), .B(n390), .Y(n304) );
  OAI221XL U1217 ( .A0(n118), .A1(n380), .B0(n119), .B1(n387), .C0(n300), .Y(
        in1[25]) );
  NAND2X1 U1218 ( .A(read_data1_out[25]), .B(n390), .Y(n300) );
  OAI221XL U1219 ( .A0(n115), .A1(n380), .B0(n116), .B1(n386), .C0(n299), .Y(
        in1[26]) );
  NAND2X1 U1220 ( .A(read_data1_out[26]), .B(n389), .Y(n299) );
  OAI221XL U1221 ( .A0(n112), .A1(n380), .B0(n113), .B1(n386), .C0(n298), .Y(
        in1[27]) );
  NAND2X1 U1222 ( .A(read_data1_out[27]), .B(n390), .Y(n298) );
  OAI221XL U1223 ( .A0(n109), .A1(n380), .B0(n110), .B1(n387), .C0(n297), .Y(
        in1[28]) );
  NAND2X1 U1224 ( .A(read_data1_out[28]), .B(n389), .Y(n297) );
  INVX1 U1225 ( .A(n430), .Y(n429) );
  INVX1 U1226 ( .A(addr2[2]), .Y(n430) );
  INVX1 U1227 ( .A(n432), .Y(n431) );
  INVX1 U1228 ( .A(addr2[3]), .Y(n432) );
  INVX1 U1229 ( .A(n426), .Y(n425) );
  INVX1 U1230 ( .A(addr2[0]), .Y(n426) );
  INVX1 U1231 ( .A(n428), .Y(n427) );
  INVX1 U1232 ( .A(addr2[1]), .Y(n428) );
  INVX1 U1233 ( .A(sel_data2_in), .Y(n211) );
  OAI2BB2X1 U1234 ( .B0(n169), .B1(n397), .A0N(read_data2[0]), .A1N(n399), .Y(
        read_data2_in[0]) );
  OAI2BB2X1 U1235 ( .B0(n136), .B1(n399), .A0N(read_data2[1]), .A1N(n399), .Y(
        read_data2_in[1]) );
  OAI2BB2X1 U1236 ( .B0(n103), .B1(n399), .A0N(read_data2[2]), .A1N(n399), .Y(
        read_data2_in[2]) );
  OAI2BB2X1 U1237 ( .B0(n94), .B1(n398), .A0N(read_data2[3]), .A1N(n399), .Y(
        read_data2_in[3]) );
  OAI2BB2X1 U1238 ( .B0(n91), .B1(n398), .A0N(read_data2[4]), .A1N(n398), .Y(
        read_data2_in[4]) );
  OAI2BB2X1 U1239 ( .B0(n88), .B1(n397), .A0N(read_data2[5]), .A1N(n398), .Y(
        read_data2_in[5]) );
  OAI2BB2X1 U1240 ( .B0(n85), .B1(n399), .A0N(read_data2[6]), .A1N(n398), .Y(
        read_data2_in[6]) );
  OAI2BB2X1 U1241 ( .B0(n82), .B1(n398), .A0N(read_data2[7]), .A1N(n399), .Y(
        read_data2_in[7]) );
  OAI2BB2X1 U1242 ( .B0(n79), .B1(n399), .A0N(read_data2[8]), .A1N(n399), .Y(
        read_data2_in[8]) );
  OAI2BB2X1 U1243 ( .B0(n73), .B1(n399), .A0N(read_data2[9]), .A1N(n398), .Y(
        read_data2_in[9]) );
  OAI2BB2X1 U1244 ( .B0(n166), .B1(n397), .A0N(read_data2[10]), .A1N(n399), 
        .Y(read_data2_in[10]) );
  OAI2BB2X1 U1245 ( .B0(n163), .B1(n398), .A0N(read_data2[11]), .A1N(n398), 
        .Y(read_data2_in[11]) );
  OAI2BB2X1 U1246 ( .B0(n160), .B1(n397), .A0N(read_data2[12]), .A1N(n398), 
        .Y(read_data2_in[12]) );
  OAI2BB2X1 U1247 ( .B0(n157), .B1(n398), .A0N(read_data2[13]), .A1N(n399), 
        .Y(read_data2_in[13]) );
  OAI2BB2X1 U1248 ( .B0(n154), .B1(n399), .A0N(read_data2[14]), .A1N(n398), 
        .Y(read_data2_in[14]) );
  OAI2BB2X1 U1249 ( .B0(n151), .B1(n397), .A0N(read_data2[15]), .A1N(n399), 
        .Y(read_data2_in[15]) );
  OAI2BB2X1 U1250 ( .B0(n148), .B1(n397), .A0N(read_data2[16]), .A1N(n399), 
        .Y(read_data2_in[16]) );
  OAI2BB2X1 U1251 ( .B0(n145), .B1(n398), .A0N(read_data2[17]), .A1N(n398), 
        .Y(read_data2_in[17]) );
  OAI2BB2X1 U1252 ( .B0(n142), .B1(n399), .A0N(read_data2[18]), .A1N(n398), 
        .Y(read_data2_in[18]) );
  OAI2BB2X1 U1253 ( .B0(n139), .B1(n397), .A0N(read_data2[19]), .A1N(n399), 
        .Y(read_data2_in[19]) );
  OAI2BB2X1 U1254 ( .B0(n133), .B1(n397), .A0N(read_data2[20]), .A1N(n398), 
        .Y(read_data2_in[20]) );
  OAI2BB2X1 U1255 ( .B0(n130), .B1(n398), .A0N(read_data2[21]), .A1N(n399), 
        .Y(read_data2_in[21]) );
  OAI2BB2X1 U1256 ( .B0(n127), .B1(n397), .A0N(read_data2[22]), .A1N(n398), 
        .Y(read_data2_in[22]) );
  OAI2BB2X1 U1257 ( .B0(n124), .B1(n398), .A0N(read_data2[23]), .A1N(n398), 
        .Y(read_data2_in[23]) );
  OAI2BB2X1 U1258 ( .B0(n121), .B1(n398), .A0N(read_data2[24]), .A1N(n398), 
        .Y(read_data2_in[24]) );
  OAI2BB2X1 U1259 ( .B0(n118), .B1(n397), .A0N(read_data2[25]), .A1N(n399), 
        .Y(read_data2_in[25]) );
  OAI2BB2X1 U1260 ( .B0(n115), .B1(n397), .A0N(read_data2[26]), .A1N(n398), 
        .Y(read_data2_in[26]) );
  OAI2BB2X1 U1261 ( .B0(n112), .B1(n397), .A0N(read_data2[27]), .A1N(n398), 
        .Y(read_data2_in[27]) );
  OAI2BB2X1 U1262 ( .B0(n109), .B1(n397), .A0N(read_data2[28]), .A1N(n399), 
        .Y(read_data2_in[28]) );
  OAI2BB2X1 U1263 ( .B0(n106), .B1(n397), .A0N(read_data2[29]), .A1N(n398), 
        .Y(read_data2_in[29]) );
  OAI2BB2X1 U1264 ( .B0(n100), .B1(n397), .A0N(read_data2[30]), .A1N(n399), 
        .Y(read_data2_in[30]) );
  OAI2BB2X1 U1265 ( .B0(n97), .B1(n399), .A0N(read_data2[31]), .A1N(n399), .Y(
        read_data2_in[31]) );
  NOR2BX1 U1266 ( .AN(funct_in_control[2]), .B(stall), .Y(funct_in[2]) );
  NOR2BX1 U1267 ( .AN(funct_in_control[3]), .B(stall), .Y(funct_in[3]) );
  INVX1 U1268 ( .A(N33), .Y(n72) );
  INVX1 U1269 ( .A(rst), .Y(N33) );
  INVX1 U1270 ( .A(n400), .Y(n403) );
  INVX1 U1271 ( .A(n400), .Y(n404) );
  INVX1 U1272 ( .A(n401), .Y(n405) );
  INVX1 U1273 ( .A(n401), .Y(n406) );
  INVX1 U1274 ( .A(n402), .Y(n407) );
endmodule

